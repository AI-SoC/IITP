module picorv32_regs(
  output rdata1[0]
  output rdata1[1]
  output rdata1[2]
  output rdata1[3]
  output rdata1[4]
  output rdata1[5]
  output rdata1[6]
  output rdata1[7]
  output rdata1[8]
  output rdata1[9]
  output rdata1[10]
  output rdata1[11]
  output rdata1[12]
  output rdata1[13]
  output rdata1[14]
  output rdata1[15]
  output rdata1[16]
  output rdata1[17]
  output rdata1[18]
  output rdata1[19]
  output rdata1[20]
  output rdata1[21]
  output rdata1[22]
  output rdata1[23]
  output rdata1[24]
  output rdata1[25]
  output rdata1[26]
  output rdata1[27]
  output rdata1[28]
  output rdata1[29]
  output rdata1[30]
  output rdata1[31]
  output rdata2[0]
  output rdata2[1]
  output rdata2[2]
  output rdata2[3]
  output rdata2[4]
  output rdata2[5]
  output rdata2[6]
  output rdata2[7]
  output rdata2[8]
  output rdata2[9]
  output rdata2[10]
  output rdata2[11]
  output rdata2[12]
  output rdata2[13]
  output rdata2[14]
  output rdata2[15]
  output rdata2[16]
  output rdata2[17]
  output rdata2[18]
  output rdata2[19]
  output rdata2[20]
  output rdata2[21]
  output rdata2[22]
  output rdata2[23]
  output rdata2[24]
  output rdata2[25]
  output rdata2[26]
  output rdata2[27]
  output rdata2[28]
  output rdata2[29]
  output rdata2[30]
  output rdata2[31]
);
  BUFX4 BUFX4_1 (.gnd(gnd), .A(raddr2_1_bF_buf14_), .Y(raddr2_1_bF_buf14_bF_buf3_), .vdd(vdd), );
  BUFX4 BUFX4_2 (.Y(raddr2_1_bF_buf14_bF_buf2_), .A(raddr2_1_bF_buf14_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_3 (.gnd(gnd), .A(raddr2_1_bF_buf14_), .Y(raddr2_1_bF_buf14_bF_buf1_), .vdd(vdd), );
  BUFX4 BUFX4_4 (.Y(raddr2_1_bF_buf14_bF_buf0_), .A(raddr2_1_bF_buf14_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_5 (.gnd(gnd), .A(clk), .Y(clk_hier0_bF_buf8), .vdd(vdd), );
  BUFX4 BUFX4_6 (.gnd(gnd), .A(clk), .Y(clk_hier0_bF_buf7), .vdd(vdd), );
  BUFX4 BUFX4_7 (.Y(clk_hier0_bF_buf6), .A(clk), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_8 (.Y(clk_hier0_bF_buf5), .A(clk), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_9 (.Y(clk_hier0_bF_buf4), .A(clk), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_10 (.gnd(gnd), .A(clk), .Y(clk_hier0_bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_11 (.gnd(gnd), .A(clk), .Y(clk_hier0_bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_12 (.gnd(gnd), .A(clk), .Y(clk_hier0_bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_13 (.gnd(gnd), .A(clk), .Y(clk_hier0_bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_14 (.Y(raddr1_1_bF_buf13_bF_buf3_), .A(raddr1_1_bF_buf13_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_15 (.Y(raddr1_1_bF_buf13_bF_buf2_), .A(raddr1_1_bF_buf13_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_16 (.Y(raddr1_1_bF_buf13_bF_buf1_), .A(raddr1_1_bF_buf13_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_17 (.Y(raddr1_1_bF_buf13_bF_buf0_), .A(raddr1_1_bF_buf13_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_18 (.Y(raddr1_1_bF_buf10_bF_buf3_), .A(raddr1_1_bF_buf10_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_19 (.Y(raddr1_1_bF_buf10_bF_buf2_), .A(raddr1_1_bF_buf10_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_20 (.gnd(gnd), .A(raddr1_1_bF_buf10_), .Y(raddr1_1_bF_buf10_bF_buf1_), .vdd(vdd), );
  BUFX4 BUFX4_21 (.gnd(gnd), .A(raddr1_1_bF_buf10_), .Y(raddr1_1_bF_buf10_bF_buf0_), .vdd(vdd), );
  BUFX4 BUFX4_22 (.gnd(gnd), .A(raddr2[0]), .Y(raddr2_0__hier0_bF_buf8), .vdd(vdd), );
  BUFX4 BUFX4_23 (.gnd(gnd), .A(raddr2[0]), .Y(raddr2_0__hier0_bF_buf7), .vdd(vdd), );
  BUFX4 BUFX4_24 (.gnd(gnd), .A(raddr2[0]), .Y(raddr2_0__hier0_bF_buf6), .vdd(vdd), );
  BUFX4 BUFX4_25 (.gnd(gnd), .A(raddr2[0]), .Y(raddr2_0__hier0_bF_buf5), .vdd(vdd), );
  BUFX4 BUFX4_26 (.gnd(gnd), .A(raddr2[0]), .Y(raddr2_0__hier0_bF_buf4), .vdd(vdd), );
  BUFX4 BUFX4_27 (.gnd(gnd), .A(raddr2[0]), .Y(raddr2_0__hier0_bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_28 (.gnd(gnd), .A(raddr2[0]), .Y(raddr2_0__hier0_bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_29 (.Y(raddr2_0__hier0_bF_buf1), .A(raddr2[0]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_30 (.Y(raddr2_0__hier0_bF_buf0), .A(raddr2[0]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_31 (.Y(raddr1_1_bF_buf9_bF_buf3_), .A(raddr1_1_bF_buf9_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_32 (.Y(raddr1_1_bF_buf9_bF_buf2_), .A(raddr1_1_bF_buf9_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_33 (.Y(raddr1_1_bF_buf9_bF_buf1_), .A(raddr1_1_bF_buf9_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_34 (.Y(raddr1_1_bF_buf9_bF_buf0_), .A(raddr1_1_bF_buf9_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_35 (.Y(raddr1_0__hier0_bF_buf8), .A(raddr1[0]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_36 (.Y(raddr1_0__hier0_bF_buf7), .A(raddr1[0]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_37 (.Y(raddr1_0__hier0_bF_buf6), .A(raddr1[0]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_38 (.Y(raddr1_0__hier0_bF_buf5), .A(raddr1[0]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_39 (.Y(raddr1_0__hier0_bF_buf4), .A(raddr1[0]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_40 (.Y(raddr1_0__hier0_bF_buf3), .A(raddr1[0]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_41 (.Y(raddr1_0__hier0_bF_buf2), .A(raddr1[0]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_42 (.Y(raddr1_0__hier0_bF_buf1), .A(raddr1[0]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_43 (.gnd(gnd), .A(raddr1[0]), .Y(raddr1_0__hier0_bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_44 (.gnd(gnd), .A(raddr2_1_bF_buf13_), .Y(raddr2_1_bF_buf13_bF_buf3_), .vdd(vdd), );
  BUFX4 BUFX4_45 (.gnd(gnd), .A(raddr2_1_bF_buf13_), .Y(raddr2_1_bF_buf13_bF_buf2_), .vdd(vdd), );
  BUFX4 BUFX4_46 (.gnd(gnd), .A(raddr2_1_bF_buf13_), .Y(raddr2_1_bF_buf13_bF_buf1_), .vdd(vdd), );
  BUFX4 BUFX4_47 (.gnd(gnd), .A(raddr2_1_bF_buf13_), .Y(raddr2_1_bF_buf13_bF_buf0_), .vdd(vdd), );
  BUFX4 BUFX4_48 (.gnd(gnd), .A(raddr1_1_bF_buf12_), .Y(raddr1_1_bF_buf12_bF_buf3_), .vdd(vdd), );
  BUFX4 BUFX4_49 (.gnd(gnd), .A(raddr1_1_bF_buf12_), .Y(raddr1_1_bF_buf12_bF_buf2_), .vdd(vdd), );
  BUFX4 BUFX4_50 (.gnd(gnd), .A(raddr1_1_bF_buf12_), .Y(raddr1_1_bF_buf12_bF_buf1_), .vdd(vdd), );
  BUFX4 BUFX4_51 (.gnd(gnd), .A(raddr1_1_bF_buf12_), .Y(raddr1_1_bF_buf12_bF_buf0_), .vdd(vdd), );
  BUFX4 BUFX4_52 (.gnd(gnd), .A(raddr2_1_bF_buf12_), .Y(raddr2_1_bF_buf12_bF_buf3_), .vdd(vdd), );
  BUFX4 BUFX4_53 (.gnd(gnd), .A(raddr2_1_bF_buf12_), .Y(raddr2_1_bF_buf12_bF_buf2_), .vdd(vdd), );
  BUFX4 BUFX4_54 (.gnd(gnd), .A(raddr2_1_bF_buf12_), .Y(raddr2_1_bF_buf12_bF_buf1_), .vdd(vdd), );
  BUFX4 BUFX4_55 (.gnd(gnd), .A(raddr2_1_bF_buf12_), .Y(raddr2_1_bF_buf12_bF_buf0_), .vdd(vdd), );
  BUFX4 BUFX4_56 (.gnd(gnd), .A(raddr1_1_bF_buf14_), .Y(raddr1_1_bF_buf14_bF_buf3_), .vdd(vdd), );
  BUFX4 BUFX4_57 (.gnd(gnd), .A(raddr1_1_bF_buf14_), .Y(raddr1_1_bF_buf14_bF_buf2_), .vdd(vdd), );
  BUFX4 BUFX4_58 (.gnd(gnd), .A(raddr1_1_bF_buf14_), .Y(raddr1_1_bF_buf14_bF_buf1_), .vdd(vdd), );
  BUFX4 BUFX4_59 (.gnd(gnd), .A(raddr1_1_bF_buf14_), .Y(raddr1_1_bF_buf14_bF_buf0_), .vdd(vdd), );
  BUFX4 BUFX4_60 (.gnd(gnd), .A(raddr1_1_bF_buf11_), .Y(raddr1_1_bF_buf11_bF_buf3_), .vdd(vdd), );
  BUFX4 BUFX4_61 (.gnd(gnd), .A(raddr1_1_bF_buf11_), .Y(raddr1_1_bF_buf11_bF_buf2_), .vdd(vdd), );
  BUFX4 BUFX4_62 (.gnd(gnd), .A(raddr1_1_bF_buf11_), .Y(raddr1_1_bF_buf11_bF_buf1_), .vdd(vdd), );
  BUFX4 BUFX4_63 (.gnd(gnd), .A(raddr1_1_bF_buf11_), .Y(raddr1_1_bF_buf11_bF_buf0_), .vdd(vdd), );
  BUFX4 BUFX4_64 (.Y(_2101__bF_buf7), .A(_2101_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_65 (.Y(_2101__bF_buf6), .A(_2101_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_66 (.Y(_2101__bF_buf5), .A(_2101_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_67 (.Y(_2101__bF_buf4), .A(_2101_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_68 (.Y(_2101__bF_buf3), .A(_2101_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_69 (.Y(_2101__bF_buf2), .A(_2101_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_70 (.Y(_2101__bF_buf1), .A(_2101_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_71 (.Y(_2101__bF_buf0), .A(_2101_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_72 (.Y(_2365__bF_buf4), .A(_2365_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_73 (.Y(_2365__bF_buf3), .A(_2365_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_74 (.Y(_2365__bF_buf2), .A(_2365_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_75 (.Y(_2365__bF_buf1), .A(_2365_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_76 (.Y(_2365__bF_buf0), .A(_2365_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_77 (.Y(_1025__bF_buf3), .A(_1025_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_78 (.Y(_1025__bF_buf2), .A(_1025_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_79 (.Y(_1025__bF_buf1), .A(_1025_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_80 (.Y(_1025__bF_buf0), .A(_1025_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_81 (.Y(raddr2_4_bF_buf4_), .A(raddr2[4]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_82 (.Y(raddr2_4_bF_buf3_), .A(raddr2[4]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_83 (.Y(raddr2_4_bF_buf2_), .A(raddr2[4]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_84 (.Y(raddr2_4_bF_buf1_), .A(raddr2[4]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_85 (.Y(raddr2_4_bF_buf0_), .A(raddr2[4]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_86 (.Y(_1063__bF_buf3), .A(_1063_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_87 (.Y(_1063__bF_buf2), .A(_1063_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_88 (.Y(_1063__bF_buf1), .A(_1063_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_89 (.Y(_1063__bF_buf0), .A(_1063_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_90 (.Y(_1310__bF_buf7), .A(_1310_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_91 (.Y(_1310__bF_buf6), .A(_1310_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_92 (.Y(_1310__bF_buf5), .A(_1310_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_93 (.Y(_1310__bF_buf4), .A(_1310_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_94 (.Y(_1310__bF_buf3), .A(_1310_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_95 (.gnd(gnd), .A(_1310_), .Y(_1310__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_96 (.gnd(gnd), .A(_1310_), .Y(_1310__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_97 (.gnd(gnd), .A(_1310_), .Y(_1310__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_98 (.gnd(gnd), .A(raddr2[1]), .Y(raddr2_1_bF_buf14_), .vdd(vdd), );
  BUFX4 BUFX4_99 (.gnd(gnd), .A(raddr2[1]), .Y(raddr2_1_bF_buf13_), .vdd(vdd), );
  BUFX4 BUFX4_100 (.gnd(gnd), .A(raddr2[1]), .Y(raddr2_1_bF_buf12_), .vdd(vdd), );
  BUFX4 BUFX4_101 (.gnd(gnd), .A(raddr2[1]), .Y(raddr2_1_bF_buf11_), .vdd(vdd), );
  BUFX4 BUFX4_102 (.gnd(gnd), .A(raddr2[1]), .Y(raddr2_1_bF_buf10_), .vdd(vdd), );
  BUFX4 BUFX4_103 (.gnd(gnd), .A(raddr2[1]), .Y(raddr2_1_bF_buf9_), .vdd(vdd), );
  BUFX4 BUFX4_104 (.gnd(gnd), .A(raddr2[1]), .Y(raddr2_1_bF_buf8_), .vdd(vdd), );
  BUFX4 BUFX4_105 (.gnd(gnd), .A(raddr2[1]), .Y(raddr2_1_bF_buf7_), .vdd(vdd), );
  BUFX4 BUFX4_106 (.gnd(gnd), .A(raddr2[1]), .Y(raddr2_1_bF_buf6_), .vdd(vdd), );
  BUFX4 BUFX4_107 (.gnd(gnd), .A(raddr2[1]), .Y(raddr2_1_bF_buf5_), .vdd(vdd), );
  BUFX4 BUFX4_108 (.gnd(gnd), .A(raddr2[1]), .Y(raddr2_1_bF_buf4_), .vdd(vdd), );
  BUFX4 BUFX4_109 (.gnd(gnd), .A(raddr2[1]), .Y(raddr2_1_bF_buf3_), .vdd(vdd), );
  BUFX4 BUFX4_110 (.gnd(gnd), .A(raddr2[1]), .Y(raddr2_1_bF_buf2_), .vdd(vdd), );
  BUFX4 BUFX4_111 (.gnd(gnd), .A(raddr2[1]), .Y(raddr2_1_bF_buf1_), .vdd(vdd), );
  BUFX4 BUFX4_112 (.gnd(gnd), .A(raddr2[1]), .Y(raddr2_1_bF_buf0_), .vdd(vdd), );
  BUFX4 BUFX4_113 (.gnd(gnd), .A(_2265_), .Y(_2265__bF_buf4), .vdd(vdd), );
  BUFX4 BUFX4_114 (.gnd(gnd), .A(_2265_), .Y(_2265__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_115 (.gnd(gnd), .A(_2265_), .Y(_2265__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_116 (.gnd(gnd), .A(_2265_), .Y(_2265__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_117 (.gnd(gnd), .A(_2265_), .Y(_2265__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_118 (.gnd(gnd), .A(raddr1[4]), .Y(raddr1_4_bF_buf4_), .vdd(vdd), );
  BUFX4 BUFX4_119 (.gnd(gnd), .A(raddr1[4]), .Y(raddr1_4_bF_buf3_), .vdd(vdd), );
  BUFX4 BUFX4_120 (.gnd(gnd), .A(raddr1[4]), .Y(raddr1_4_bF_buf2_), .vdd(vdd), );
  BUFX4 BUFX4_121 (.gnd(gnd), .A(raddr1[4]), .Y(raddr1_4_bF_buf1_), .vdd(vdd), );
  BUFX4 BUFX4_122 (.gnd(gnd), .A(raddr1[4]), .Y(raddr1_4_bF_buf0_), .vdd(vdd), );
  BUFX4 BUFX4_123 (.gnd(gnd), .A(_1019_), .Y(_1019__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_124 (.gnd(gnd), .A(_1019_), .Y(_1019__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_125 (.gnd(gnd), .A(_1019_), .Y(_1019__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_126 (.gnd(gnd), .A(_1019_), .Y(_1019__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_127 (.gnd(gnd), .A(_999_), .Y(_999__bF_buf4), .vdd(vdd), );
  BUFX4 BUFX4_128 (.gnd(gnd), .A(_999_), .Y(_999__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_129 (.gnd(gnd), .A(_999_), .Y(_999__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_130 (.gnd(gnd), .A(_999_), .Y(_999__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_131 (.gnd(gnd), .A(_999_), .Y(_999__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_132 (.gnd(gnd), .A(_1057_), .Y(_1057__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_133 (.gnd(gnd), .A(_1057_), .Y(_1057__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_134 (.gnd(gnd), .A(_1057_), .Y(_1057__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_135 (.gnd(gnd), .A(_1057_), .Y(_1057__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_136 (.gnd(gnd), .A(_2415_), .Y(_2415__bF_buf8), .vdd(vdd), );
  BUFX4 BUFX4_137 (.gnd(gnd), .A(_2415_), .Y(_2415__bF_buf7), .vdd(vdd), );
  BUFX4 BUFX4_138 (.gnd(gnd), .A(_2415_), .Y(_2415__bF_buf6), .vdd(vdd), );
  BUFX4 BUFX4_139 (.gnd(gnd), .A(_2415_), .Y(_2415__bF_buf5), .vdd(vdd), );
  BUFX4 BUFX4_140 (.gnd(gnd), .A(_2415_), .Y(_2415__bF_buf4), .vdd(vdd), );
  BUFX4 BUFX4_141 (.gnd(gnd), .A(_2415_), .Y(_2415__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_142 (.Y(_2415__bF_buf2), .A(_2415_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_143 (.Y(_2415__bF_buf1), .A(_2415_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_144 (.Y(_2415__bF_buf0), .A(_2415_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_145 (.Y(raddr1_1_bF_buf14_), .A(raddr1[1]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_146 (.Y(raddr1_1_bF_buf13_), .A(raddr1[1]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_147 (.Y(raddr1_1_bF_buf12_), .A(raddr1[1]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_148 (.Y(raddr1_1_bF_buf11_), .A(raddr1[1]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_149 (.Y(raddr1_1_bF_buf10_), .A(raddr1[1]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_150 (.Y(raddr1_1_bF_buf9_), .A(raddr1[1]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_151 (.Y(raddr1_1_bF_buf8_), .A(raddr1[1]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_152 (.Y(raddr1_1_bF_buf7_), .A(raddr1[1]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_153 (.Y(raddr1_1_bF_buf6_), .A(raddr1[1]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_154 (.Y(raddr1_1_bF_buf5_), .A(raddr1[1]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_155 (.Y(raddr1_1_bF_buf4_), .A(raddr1[1]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_156 (.Y(raddr1_1_bF_buf3_), .A(raddr1[1]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_157 (.Y(raddr1_1_bF_buf2_), .A(raddr1[1]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_158 (.Y(raddr1_1_bF_buf1_), .A(raddr1[1]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_159 (.Y(raddr1_1_bF_buf0_), .A(raddr1[1]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_160 (.Y(_1571__bF_buf7), .A(_1571_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_161 (.Y(_1571__bF_buf6), .A(_1571_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_162 (.Y(_1571__bF_buf5), .A(_1571_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_163 (.Y(_1571__bF_buf4), .A(_1571_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_164 (.Y(_1571__bF_buf3), .A(_1571_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_165 (.Y(_1571__bF_buf2), .A(_1571_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_166 (.Y(_1571__bF_buf1), .A(_1571_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_167 (.Y(_1571__bF_buf0), .A(_1571_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_168 (.Y(_1207__bF_buf7), .A(_1207_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_169 (.Y(_1207__bF_buf6), .A(_1207_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_170 (.Y(_1207__bF_buf5), .A(_1207_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_171 (.Y(_1207__bF_buf4), .A(_1207_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_172 (.Y(_1207__bF_buf3), .A(_1207_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_173 (.Y(_1207__bF_buf2), .A(_1207_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_174 (.Y(_1207__bF_buf1), .A(_1207_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_175 (.Y(_1207__bF_buf0), .A(_1207_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_176 (.Y(_2165__bF_buf4), .A(_2165_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_177 (.Y(_2165__bF_buf3), .A(_2165_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_178 (.Y(_2165__bF_buf2), .A(_2165_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_179 (.Y(_2165__bF_buf1), .A(_2165_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_180 (.Y(_2165__bF_buf0), .A(_2165_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_181 (.Y(_1013__bF_buf3), .A(_1013_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_182 (.Y(_1013__bF_buf2), .A(_1013_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_183 (.Y(_1013__bF_buf1), .A(_1013_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_184 (.Y(_1013__bF_buf0), .A(_1013_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_185 (.Y(_1051__bF_buf3), .A(_1051_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_186 (.Y(_1051__bF_buf2), .A(_1051_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_187 (.Y(_1051__bF_buf1), .A(_1051_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_188 (.Y(_1051__bF_buf0), .A(_1051_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_189 (.Y(_1374__bF_buf7), .A(_1374_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_190 (.Y(_1374__bF_buf6), .A(_1374_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_191 (.Y(_1374__bF_buf5), .A(_1374_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_192 (.Y(_1374__bF_buf4), .A(_1374_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_193 (.Y(_1374__bF_buf3), .A(_1374_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_194 (.Y(_1374__bF_buf2), .A(_1374_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_195 (.Y(_1374__bF_buf1), .A(_1374_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_196 (.Y(_1374__bF_buf0), .A(_1374_), .gnd(gnd), .vdd(vdd), );
  CLKBUF1 CLKBUF1_1 (.Y(clk_bF_buf98), .A(clk_hier0_bF_buf8), .gnd(gnd), .vdd(vdd), );
  CLKBUF1 CLKBUF1_2 (.Y(clk_bF_buf97), .A(clk_hier0_bF_buf7), .gnd(gnd), .vdd(vdd), );
  CLKBUF1 CLKBUF1_3 (.Y(clk_bF_buf96), .A(clk_hier0_bF_buf6), .gnd(gnd), .vdd(vdd), );
  CLKBUF1 CLKBUF1_4 (.Y(clk_bF_buf95), .A(clk_hier0_bF_buf5), .gnd(gnd), .vdd(vdd), );
  CLKBUF1 CLKBUF1_5 (.Y(clk_bF_buf94), .A(clk_hier0_bF_buf4), .gnd(gnd), .vdd(vdd), );
  CLKBUF1 CLKBUF1_6 (.Y(clk_bF_buf93), .A(clk_hier0_bF_buf3), .gnd(gnd), .vdd(vdd), );
  CLKBUF1 CLKBUF1_7 (.Y(clk_bF_buf92), .A(clk_hier0_bF_buf2), .gnd(gnd), .vdd(vdd), );
  CLKBUF1 CLKBUF1_8 (.Y(clk_bF_buf91), .A(clk_hier0_bF_buf1), .gnd(gnd), .vdd(vdd), );
  CLKBUF1 CLKBUF1_9 (.Y(clk_bF_buf90), .A(clk_hier0_bF_buf0), .gnd(gnd), .vdd(vdd), );
  CLKBUF1 CLKBUF1_10 (.Y(clk_bF_buf89), .A(clk_hier0_bF_buf8), .gnd(gnd), .vdd(vdd), );
  CLKBUF1 CLKBUF1_11 (.Y(clk_bF_buf88), .A(clk_hier0_bF_buf7), .gnd(gnd), .vdd(vdd), );
  CLKBUF1 CLKBUF1_12 (.Y(clk_bF_buf87), .A(clk_hier0_bF_buf6), .gnd(gnd), .vdd(vdd), );
  CLKBUF1 CLKBUF1_13 (.Y(clk_bF_buf86), .A(clk_hier0_bF_buf5), .gnd(gnd), .vdd(vdd), );
  CLKBUF1 CLKBUF1_14 (.Y(clk_bF_buf85), .A(clk_hier0_bF_buf4), .gnd(gnd), .vdd(vdd), );
  CLKBUF1 CLKBUF1_15 (.Y(clk_bF_buf84), .A(clk_hier0_bF_buf3), .gnd(gnd), .vdd(vdd), );
  CLKBUF1 CLKBUF1_16 (.gnd(gnd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf83), .vdd(vdd), );
  CLKBUF1 CLKBUF1_17 (.gnd(gnd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf82), .vdd(vdd), );
  CLKBUF1 CLKBUF1_18 (.gnd(gnd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf81), .vdd(vdd), );
  CLKBUF1 CLKBUF1_19 (.gnd(gnd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf80), .vdd(vdd), );
  CLKBUF1 CLKBUF1_20 (.gnd(gnd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf79), .vdd(vdd), );
  CLKBUF1 CLKBUF1_21 (.gnd(gnd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf78), .vdd(vdd), );
  CLKBUF1 CLKBUF1_22 (.gnd(gnd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf77), .vdd(vdd), );
  CLKBUF1 CLKBUF1_23 (.gnd(gnd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf76), .vdd(vdd), );
  CLKBUF1 CLKBUF1_24 (.gnd(gnd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf75), .vdd(vdd), );
  CLKBUF1 CLKBUF1_25 (.gnd(gnd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf74), .vdd(vdd), );
  CLKBUF1 CLKBUF1_26 (.gnd(gnd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf73), .vdd(vdd), );
  CLKBUF1 CLKBUF1_27 (.gnd(gnd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf72), .vdd(vdd), );
  CLKBUF1 CLKBUF1_28 (.gnd(gnd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf71), .vdd(vdd), );
  CLKBUF1 CLKBUF1_29 (.gnd(gnd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf70), .vdd(vdd), );
  CLKBUF1 CLKBUF1_30 (.gnd(gnd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf69), .vdd(vdd), );
  CLKBUF1 CLKBUF1_31 (.gnd(gnd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf68), .vdd(vdd), );
  CLKBUF1 CLKBUF1_32 (.gnd(gnd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf67), .vdd(vdd), );
  CLKBUF1 CLKBUF1_33 (.gnd(gnd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf66), .vdd(vdd), );
  CLKBUF1 CLKBUF1_34 (.gnd(gnd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf65), .vdd(vdd), );
  CLKBUF1 CLKBUF1_35 (.gnd(gnd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf64), .vdd(vdd), );
  CLKBUF1 CLKBUF1_36 (.gnd(gnd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf63), .vdd(vdd), );
  CLKBUF1 CLKBUF1_37 (.gnd(gnd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf62), .vdd(vdd), );
  CLKBUF1 CLKBUF1_38 (.gnd(gnd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf61), .vdd(vdd), );
  CLKBUF1 CLKBUF1_39 (.gnd(gnd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf60), .vdd(vdd), );
  CLKBUF1 CLKBUF1_40 (.gnd(gnd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf59), .vdd(vdd), );
  CLKBUF1 CLKBUF1_41 (.gnd(gnd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf58), .vdd(vdd), );
  CLKBUF1 CLKBUF1_42 (.gnd(gnd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf57), .vdd(vdd), );
  CLKBUF1 CLKBUF1_43 (.gnd(gnd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf56), .vdd(vdd), );
  CLKBUF1 CLKBUF1_44 (.gnd(gnd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf55), .vdd(vdd), );
  CLKBUF1 CLKBUF1_45 (.gnd(gnd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf54), .vdd(vdd), );
  CLKBUF1 CLKBUF1_46 (.gnd(gnd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf53), .vdd(vdd), );
  CLKBUF1 CLKBUF1_47 (.gnd(gnd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf52), .vdd(vdd), );
  CLKBUF1 CLKBUF1_48 (.gnd(gnd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf51), .vdd(vdd), );
  CLKBUF1 CLKBUF1_49 (.gnd(gnd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf50), .vdd(vdd), );
  CLKBUF1 CLKBUF1_50 (.gnd(gnd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf49), .vdd(vdd), );
  CLKBUF1 CLKBUF1_51 (.gnd(gnd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf48), .vdd(vdd), );
  CLKBUF1 CLKBUF1_52 (.gnd(gnd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf47), .vdd(vdd), );
  CLKBUF1 CLKBUF1_53 (.gnd(gnd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf46), .vdd(vdd), );
  CLKBUF1 CLKBUF1_54 (.gnd(gnd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf45), .vdd(vdd), );
  CLKBUF1 CLKBUF1_55 (.gnd(gnd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf44), .vdd(vdd), );
  CLKBUF1 CLKBUF1_56 (.gnd(gnd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf43), .vdd(vdd), );
  CLKBUF1 CLKBUF1_57 (.gnd(gnd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf42), .vdd(vdd), );
  CLKBUF1 CLKBUF1_58 (.gnd(gnd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf41), .vdd(vdd), );
  CLKBUF1 CLKBUF1_59 (.gnd(gnd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf40), .vdd(vdd), );
  CLKBUF1 CLKBUF1_60 (.gnd(gnd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf39), .vdd(vdd), );
  CLKBUF1 CLKBUF1_61 (.gnd(gnd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf38), .vdd(vdd), );
  CLKBUF1 CLKBUF1_62 (.gnd(gnd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf37), .vdd(vdd), );
  CLKBUF1 CLKBUF1_63 (.gnd(gnd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf36), .vdd(vdd), );
  CLKBUF1 CLKBUF1_64 (.gnd(gnd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf35), .vdd(vdd), );
  CLKBUF1 CLKBUF1_65 (.gnd(gnd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf34), .vdd(vdd), );
  CLKBUF1 CLKBUF1_66 (.gnd(gnd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf33), .vdd(vdd), );
  CLKBUF1 CLKBUF1_67 (.gnd(gnd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf32), .vdd(vdd), );
  CLKBUF1 CLKBUF1_68 (.gnd(gnd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf31), .vdd(vdd), );
  CLKBUF1 CLKBUF1_69 (.gnd(gnd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf30), .vdd(vdd), );
  CLKBUF1 CLKBUF1_70 (.gnd(gnd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf29), .vdd(vdd), );
  CLKBUF1 CLKBUF1_71 (.gnd(gnd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf28), .vdd(vdd), );
  CLKBUF1 CLKBUF1_72 (.gnd(gnd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf27), .vdd(vdd), );
  CLKBUF1 CLKBUF1_73 (.gnd(gnd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf26), .vdd(vdd), );
  CLKBUF1 CLKBUF1_74 (.gnd(gnd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf25), .vdd(vdd), );
  CLKBUF1 CLKBUF1_75 (.gnd(gnd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf24), .vdd(vdd), );
  CLKBUF1 CLKBUF1_76 (.gnd(gnd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf23), .vdd(vdd), );
  CLKBUF1 CLKBUF1_77 (.gnd(gnd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf22), .vdd(vdd), );
  CLKBUF1 CLKBUF1_78 (.gnd(gnd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf21), .vdd(vdd), );
  CLKBUF1 CLKBUF1_79 (.gnd(gnd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf20), .vdd(vdd), );
  CLKBUF1 CLKBUF1_80 (.gnd(gnd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf19), .vdd(vdd), );
  CLKBUF1 CLKBUF1_81 (.gnd(gnd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf18), .vdd(vdd), );
  CLKBUF1 CLKBUF1_82 (.gnd(gnd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf17), .vdd(vdd), );
  CLKBUF1 CLKBUF1_83 (.gnd(gnd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf16), .vdd(vdd), );
  CLKBUF1 CLKBUF1_84 (.gnd(gnd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf15), .vdd(vdd), );
  CLKBUF1 CLKBUF1_85 (.gnd(gnd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf14), .vdd(vdd), );
  CLKBUF1 CLKBUF1_86 (.gnd(gnd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf13), .vdd(vdd), );
  CLKBUF1 CLKBUF1_87 (.gnd(gnd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf12), .vdd(vdd), );
  CLKBUF1 CLKBUF1_88 (.gnd(gnd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf11), .vdd(vdd), );
  CLKBUF1 CLKBUF1_89 (.gnd(gnd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf10), .vdd(vdd), );
  CLKBUF1 CLKBUF1_90 (.gnd(gnd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf9), .vdd(vdd), );
  CLKBUF1 CLKBUF1_91 (.gnd(gnd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf8), .vdd(vdd), );
  CLKBUF1 CLKBUF1_92 (.gnd(gnd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf7), .vdd(vdd), );
  CLKBUF1 CLKBUF1_93 (.gnd(gnd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf6), .vdd(vdd), );
  CLKBUF1 CLKBUF1_94 (.gnd(gnd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf5), .vdd(vdd), );
  CLKBUF1 CLKBUF1_95 (.gnd(gnd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf4), .vdd(vdd), );
  CLKBUF1 CLKBUF1_96 (.gnd(gnd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf3), .vdd(vdd), );
  CLKBUF1 CLKBUF1_97 (.gnd(gnd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf2), .vdd(vdd), );
  CLKBUF1 CLKBUF1_98 (.gnd(gnd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf1), .vdd(vdd), );
  CLKBUF1 CLKBUF1_99 (.gnd(gnd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_197 (.gnd(gnd), .A(_1104_), .Y(_1104__bF_buf14), .vdd(vdd), );
  BUFX4 BUFX4_198 (.gnd(gnd), .A(_1104_), .Y(_1104__bF_buf13), .vdd(vdd), );
  BUFX4 BUFX4_199 (.gnd(gnd), .A(_1104_), .Y(_1104__bF_buf12), .vdd(vdd), );
  BUFX4 BUFX4_200 (.gnd(gnd), .A(_1104_), .Y(_1104__bF_buf11), .vdd(vdd), );
  BUFX4 BUFX4_201 (.gnd(gnd), .A(_1104_), .Y(_1104__bF_buf10), .vdd(vdd), );
  BUFX4 BUFX4_202 (.gnd(gnd), .A(_1104_), .Y(_1104__bF_buf9), .vdd(vdd), );
  BUFX4 BUFX4_203 (.gnd(gnd), .A(_1104_), .Y(_1104__bF_buf8), .vdd(vdd), );
  BUFX4 BUFX4_204 (.gnd(gnd), .A(_1104_), .Y(_1104__bF_buf7), .vdd(vdd), );
  BUFX4 BUFX4_205 (.gnd(gnd), .A(_1104_), .Y(_1104__bF_buf6), .vdd(vdd), );
  BUFX4 BUFX4_206 (.gnd(gnd), .A(_1104_), .Y(_1104__bF_buf5), .vdd(vdd), );
  BUFX4 BUFX4_207 (.gnd(gnd), .A(_1104_), .Y(_1104__bF_buf4), .vdd(vdd), );
  BUFX4 BUFX4_208 (.gnd(gnd), .A(_1104_), .Y(_1104__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_209 (.gnd(gnd), .A(_1104_), .Y(_1104__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_210 (.gnd(gnd), .A(_1104_), .Y(_1104__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_211 (.gnd(gnd), .A(_1104_), .Y(_1104__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_212 (.gnd(gnd), .A(_1142_), .Y(_1142__bF_buf5), .vdd(vdd), );
  BUFX4 BUFX4_213 (.gnd(gnd), .A(_1142_), .Y(_1142__bF_buf4), .vdd(vdd), );
  BUFX4 BUFX4_214 (.gnd(gnd), .A(_1142_), .Y(_1142__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_215 (.gnd(gnd), .A(_1142_), .Y(_1142__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_216 (.gnd(gnd), .A(_1142_), .Y(_1142__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_217 (.gnd(gnd), .A(_1142_), .Y(_1142__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_218 (.Y(_1007__bF_buf3), .A(_1007_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_219 (.Y(_1007__bF_buf2), .A(_1007_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_220 (.Y(_1007__bF_buf1), .A(_1007_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_221 (.Y(_1007__bF_buf0), .A(_1007_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_222 (.Y(_1045__bF_buf3), .A(_1045_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_223 (.Y(_1045__bF_buf2), .A(_1045_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_224 (.Y(_1045__bF_buf1), .A(_1045_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_225 (.Y(_1045__bF_buf0), .A(_1045_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_226 (.Y(_1274__bF_buf4), .A(_1274_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_227 (.Y(_1274__bF_buf3), .A(_1274_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_228 (.Y(_1274__bF_buf2), .A(_1274_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_229 (.Y(_1274__bF_buf1), .A(_1274_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_230 (.Y(_1274__bF_buf0), .A(_1274_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_231 (.Y(_1039__bF_buf3), .A(_1039_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_232 (.Y(_1039__bF_buf2), .A(_1039_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_233 (.Y(_1039__bF_buf1), .A(_1039_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_234 (.Y(_1039__bF_buf0), .A(_1039_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_235 (.Y(_1803__bF_buf7), .A(_1803_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_236 (.Y(_1803__bF_buf6), .A(_1803_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_237 (.Y(_1803__bF_buf5), .A(_1803_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_238 (.Y(_1803__bF_buf4), .A(_1803_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_239 (.Y(_1803__bF_buf3), .A(_1803_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_240 (.Y(_1803__bF_buf2), .A(_1803_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_241 (.Y(_1803__bF_buf1), .A(_1803_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_242 (.Y(_1803__bF_buf0), .A(_1803_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_243 (.Y(_1001__bF_buf9), .A(_1001_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_244 (.Y(_1001__bF_buf8), .A(_1001_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_245 (.Y(_1001__bF_buf7), .A(_1001_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_246 (.Y(_1001__bF_buf6), .A(_1001_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_247 (.Y(_1001__bF_buf5), .A(_1001_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_248 (.Y(_1001__bF_buf4), .A(_1001_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_249 (.Y(_1001__bF_buf3), .A(_1001_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_250 (.Y(_1001__bF_buf2), .A(_1001_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_251 (.Y(_1001__bF_buf1), .A(_1001_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_252 (.Y(_1001__bF_buf0), .A(_1001_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_253 (.Y(_1033__bF_buf3), .A(_1033_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_254 (.Y(_1033__bF_buf2), .A(_1033_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_255 (.Y(_1033__bF_buf1), .A(_1033_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_256 (.Y(_1033__bF_buf0), .A(_1033_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_257 (.Y(_2332__bF_buf4), .A(_2332_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_258 (.Y(_2332__bF_buf3), .A(_2332_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_259 (.Y(_2332__bF_buf2), .A(_2332_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_260 (.Y(_2332__bF_buf1), .A(_2332_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_261 (.Y(_2332__bF_buf0), .A(_2332_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_262 (.Y(_1506__bF_buf5), .A(_1506_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_263 (.Y(_1506__bF_buf4), .A(_1506_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_264 (.Y(_1506__bF_buf3), .A(_1506_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_265 (.Y(_1506__bF_buf2), .A(_1506_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_266 (.Y(_1506__bF_buf1), .A(_1506_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_267 (.Y(_1506__bF_buf0), .A(_1506_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_268 (.Y(_1867__bF_buf4), .A(_1867_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_269 (.Y(_1867__bF_buf3), .A(_1867_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_270 (.Y(_1867__bF_buf2), .A(_1867_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_271 (.Y(_1867__bF_buf1), .A(_1867_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_272 (.Y(_1867__bF_buf0), .A(_1867_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_273 (.Y(_1027__bF_buf3), .A(_1027_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_274 (.Y(_1027__bF_buf2), .A(_1027_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_275 (.Y(_1027__bF_buf1), .A(_1027_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_276 (.Y(_1027__bF_buf0), .A(_1027_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_277 (.Y(_2100__bF_buf8), .A(_2100_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_278 (.Y(_2100__bF_buf7), .A(_2100_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_279 (.Y(_2100__bF_buf6), .A(_2100_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_280 (.Y(_2100__bF_buf5), .A(_2100_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_281 (.Y(_2100__bF_buf4), .A(_2100_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_282 (.Y(_2100__bF_buf3), .A(_2100_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_283 (.Y(_2100__bF_buf2), .A(_2100_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_284 (.Y(_2100__bF_buf1), .A(_2100_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_285 (.Y(_2100__bF_buf0), .A(_2100_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_286 (.Y(_1309__bF_buf5), .A(_1309_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_287 (.Y(_1309__bF_buf4), .A(_1309_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_288 (.Y(_1309__bF_buf3), .A(_1309_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_289 (.Y(_1309__bF_buf2), .A(_1309_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_290 (.Y(_1309__bF_buf1), .A(_1309_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_291 (.Y(_1309__bF_buf0), .A(_1309_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_292 (.Y(_2399__bF_buf8), .A(_2399_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_293 (.Y(_2399__bF_buf7), .A(_2399_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_294 (.Y(_2399__bF_buf6), .A(_2399_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_295 (.Y(_2399__bF_buf5), .A(_2399_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_296 (.Y(_2399__bF_buf4), .A(_2399_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_297 (.Y(_2399__bF_buf3), .A(_2399_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_298 (.Y(_2399__bF_buf2), .A(_2399_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_299 (.Y(_2399__bF_buf1), .A(_2399_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_300 (.Y(_2399__bF_buf0), .A(_2399_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_301 (.Y(_1059__bF_buf3), .A(_1059_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_302 (.Y(_1059__bF_buf2), .A(_1059_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_303 (.Y(_1059__bF_buf1), .A(_1059_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_304 (.Y(_1059__bF_buf0), .A(_1059_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_305 (.Y(_2000__bF_buf7), .A(_2000_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_306 (.Y(_2000__bF_buf6), .A(_2000_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_307 (.Y(_2000__bF_buf5), .A(_2000_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_308 (.Y(_2000__bF_buf4), .A(_2000_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_309 (.Y(_2000__bF_buf3), .A(_2000_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_310 (.Y(_2000__bF_buf2), .A(_2000_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_311 (.Y(_2000__bF_buf1), .A(_2000_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_312 (.Y(_2000__bF_buf0), .A(_2000_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_313 (.Y(_1021__bF_buf3), .A(_1021_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_314 (.Y(_1021__bF_buf2), .A(_1021_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_315 (.Y(_1021__bF_buf1), .A(_1021_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_316 (.Y(_1021__bF_buf0), .A(_1021_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_317 (.Y(raddr2_0_bF_buf96_), .A(raddr2_0__hier0_bF_buf8), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_318 (.Y(raddr2_0_bF_buf95_), .A(raddr2_0__hier0_bF_buf7), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_319 (.Y(raddr2_0_bF_buf94_), .A(raddr2_0__hier0_bF_buf6), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_320 (.Y(raddr2_0_bF_buf93_), .A(raddr2_0__hier0_bF_buf5), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_321 (.Y(raddr2_0_bF_buf92_), .A(raddr2_0__hier0_bF_buf4), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_322 (.Y(raddr2_0_bF_buf91_), .A(raddr2_0__hier0_bF_buf3), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_323 (.Y(raddr2_0_bF_buf90_), .A(raddr2_0__hier0_bF_buf2), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_324 (.Y(raddr2_0_bF_buf89_), .A(raddr2_0__hier0_bF_buf1), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_325 (.Y(raddr2_0_bF_buf88_), .A(raddr2_0__hier0_bF_buf0), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_326 (.Y(raddr2_0_bF_buf87_), .A(raddr2_0__hier0_bF_buf8), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_327 (.Y(raddr2_0_bF_buf86_), .A(raddr2_0__hier0_bF_buf7), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_328 (.Y(raddr2_0_bF_buf85_), .A(raddr2_0__hier0_bF_buf6), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_329 (.Y(raddr2_0_bF_buf84_), .A(raddr2_0__hier0_bF_buf5), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_330 (.Y(raddr2_0_bF_buf83_), .A(raddr2_0__hier0_bF_buf4), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_331 (.Y(raddr2_0_bF_buf82_), .A(raddr2_0__hier0_bF_buf3), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_332 (.Y(raddr2_0_bF_buf81_), .A(raddr2_0__hier0_bF_buf2), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_333 (.Y(raddr2_0_bF_buf80_), .A(raddr2_0__hier0_bF_buf1), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_334 (.Y(raddr2_0_bF_buf79_), .A(raddr2_0__hier0_bF_buf0), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_335 (.Y(raddr2_0_bF_buf78_), .A(raddr2_0__hier0_bF_buf8), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_336 (.Y(raddr2_0_bF_buf77_), .A(raddr2_0__hier0_bF_buf7), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_337 (.Y(raddr2_0_bF_buf76_), .A(raddr2_0__hier0_bF_buf6), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_338 (.Y(raddr2_0_bF_buf75_), .A(raddr2_0__hier0_bF_buf5), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_339 (.Y(raddr2_0_bF_buf74_), .A(raddr2_0__hier0_bF_buf4), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_340 (.Y(raddr2_0_bF_buf73_), .A(raddr2_0__hier0_bF_buf3), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_341 (.Y(raddr2_0_bF_buf72_), .A(raddr2_0__hier0_bF_buf2), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_342 (.Y(raddr2_0_bF_buf71_), .A(raddr2_0__hier0_bF_buf1), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_343 (.Y(raddr2_0_bF_buf70_), .A(raddr2_0__hier0_bF_buf0), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_344 (.Y(raddr2_0_bF_buf69_), .A(raddr2_0__hier0_bF_buf8), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_345 (.Y(raddr2_0_bF_buf68_), .A(raddr2_0__hier0_bF_buf7), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_346 (.Y(raddr2_0_bF_buf67_), .A(raddr2_0__hier0_bF_buf6), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_347 (.Y(raddr2_0_bF_buf66_), .A(raddr2_0__hier0_bF_buf5), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_348 (.Y(raddr2_0_bF_buf65_), .A(raddr2_0__hier0_bF_buf4), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_349 (.Y(raddr2_0_bF_buf64_), .A(raddr2_0__hier0_bF_buf3), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_350 (.Y(raddr2_0_bF_buf63_), .A(raddr2_0__hier0_bF_buf2), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_351 (.Y(raddr2_0_bF_buf62_), .A(raddr2_0__hier0_bF_buf1), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_352 (.Y(raddr2_0_bF_buf61_), .A(raddr2_0__hier0_bF_buf0), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_353 (.Y(raddr2_0_bF_buf60_), .A(raddr2_0__hier0_bF_buf8), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_354 (.Y(raddr2_0_bF_buf59_), .A(raddr2_0__hier0_bF_buf7), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_355 (.Y(raddr2_0_bF_buf58_), .A(raddr2_0__hier0_bF_buf6), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_356 (.Y(raddr2_0_bF_buf57_), .A(raddr2_0__hier0_bF_buf5), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_357 (.Y(raddr2_0_bF_buf56_), .A(raddr2_0__hier0_bF_buf4), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_358 (.Y(raddr2_0_bF_buf55_), .A(raddr2_0__hier0_bF_buf3), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_359 (.Y(raddr2_0_bF_buf54_), .A(raddr2_0__hier0_bF_buf2), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_360 (.Y(raddr2_0_bF_buf53_), .A(raddr2_0__hier0_bF_buf1), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_361 (.Y(raddr2_0_bF_buf52_), .A(raddr2_0__hier0_bF_buf0), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_362 (.Y(raddr2_0_bF_buf51_), .A(raddr2_0__hier0_bF_buf8), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_363 (.Y(raddr2_0_bF_buf50_), .A(raddr2_0__hier0_bF_buf7), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_364 (.Y(raddr2_0_bF_buf49_), .A(raddr2_0__hier0_bF_buf6), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_365 (.Y(raddr2_0_bF_buf48_), .A(raddr2_0__hier0_bF_buf5), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_366 (.Y(raddr2_0_bF_buf47_), .A(raddr2_0__hier0_bF_buf4), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_367 (.Y(raddr2_0_bF_buf46_), .A(raddr2_0__hier0_bF_buf3), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_368 (.Y(raddr2_0_bF_buf45_), .A(raddr2_0__hier0_bF_buf2), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_369 (.Y(raddr2_0_bF_buf44_), .A(raddr2_0__hier0_bF_buf1), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_370 (.Y(raddr2_0_bF_buf43_), .A(raddr2_0__hier0_bF_buf0), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_371 (.Y(raddr2_0_bF_buf42_), .A(raddr2_0__hier0_bF_buf8), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_372 (.Y(raddr2_0_bF_buf41_), .A(raddr2_0__hier0_bF_buf7), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_373 (.Y(raddr2_0_bF_buf40_), .A(raddr2_0__hier0_bF_buf6), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_374 (.Y(raddr2_0_bF_buf39_), .A(raddr2_0__hier0_bF_buf5), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_375 (.Y(raddr2_0_bF_buf38_), .A(raddr2_0__hier0_bF_buf4), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_376 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf3), .Y(raddr2_0_bF_buf37_), .vdd(vdd), );
  BUFX4 BUFX4_377 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf2), .Y(raddr2_0_bF_buf36_), .vdd(vdd), );
  BUFX4 BUFX4_378 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf1), .Y(raddr2_0_bF_buf35_), .vdd(vdd), );
  BUFX4 BUFX4_379 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf0), .Y(raddr2_0_bF_buf34_), .vdd(vdd), );
  BUFX4 BUFX4_380 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf8), .Y(raddr2_0_bF_buf33_), .vdd(vdd), );
  BUFX4 BUFX4_381 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf7), .Y(raddr2_0_bF_buf32_), .vdd(vdd), );
  BUFX4 BUFX4_382 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf6), .Y(raddr2_0_bF_buf31_), .vdd(vdd), );
  BUFX4 BUFX4_383 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf5), .Y(raddr2_0_bF_buf30_), .vdd(vdd), );
  BUFX4 BUFX4_384 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf4), .Y(raddr2_0_bF_buf29_), .vdd(vdd), );
  BUFX4 BUFX4_385 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf3), .Y(raddr2_0_bF_buf28_), .vdd(vdd), );
  BUFX4 BUFX4_386 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf2), .Y(raddr2_0_bF_buf27_), .vdd(vdd), );
  BUFX4 BUFX4_387 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf1), .Y(raddr2_0_bF_buf26_), .vdd(vdd), );
  BUFX4 BUFX4_388 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf0), .Y(raddr2_0_bF_buf25_), .vdd(vdd), );
  BUFX4 BUFX4_389 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf8), .Y(raddr2_0_bF_buf24_), .vdd(vdd), );
  BUFX4 BUFX4_390 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf7), .Y(raddr2_0_bF_buf23_), .vdd(vdd), );
  BUFX4 BUFX4_391 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf6), .Y(raddr2_0_bF_buf22_), .vdd(vdd), );
  BUFX4 BUFX4_392 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf5), .Y(raddr2_0_bF_buf21_), .vdd(vdd), );
  BUFX4 BUFX4_393 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf4), .Y(raddr2_0_bF_buf20_), .vdd(vdd), );
  BUFX4 BUFX4_394 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf3), .Y(raddr2_0_bF_buf19_), .vdd(vdd), );
  BUFX4 BUFX4_395 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf2), .Y(raddr2_0_bF_buf18_), .vdd(vdd), );
  BUFX4 BUFX4_396 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf1), .Y(raddr2_0_bF_buf17_), .vdd(vdd), );
  BUFX4 BUFX4_397 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf0), .Y(raddr2_0_bF_buf16_), .vdd(vdd), );
  BUFX4 BUFX4_398 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf8), .Y(raddr2_0_bF_buf15_), .vdd(vdd), );
  BUFX4 BUFX4_399 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf7), .Y(raddr2_0_bF_buf14_), .vdd(vdd), );
  BUFX4 BUFX4_400 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf6), .Y(raddr2_0_bF_buf13_), .vdd(vdd), );
  BUFX4 BUFX4_401 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf5), .Y(raddr2_0_bF_buf12_), .vdd(vdd), );
  BUFX4 BUFX4_402 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf4), .Y(raddr2_0_bF_buf11_), .vdd(vdd), );
  BUFX4 BUFX4_403 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf3), .Y(raddr2_0_bF_buf10_), .vdd(vdd), );
  BUFX4 BUFX4_404 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf2), .Y(raddr2_0_bF_buf9_), .vdd(vdd), );
  BUFX4 BUFX4_405 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf1), .Y(raddr2_0_bF_buf8_), .vdd(vdd), );
  BUFX4 BUFX4_406 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf0), .Y(raddr2_0_bF_buf7_), .vdd(vdd), );
  BUFX4 BUFX4_407 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf8), .Y(raddr2_0_bF_buf6_), .vdd(vdd), );
  BUFX4 BUFX4_408 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf7), .Y(raddr2_0_bF_buf5_), .vdd(vdd), );
  BUFX4 BUFX4_409 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf6), .Y(raddr2_0_bF_buf4_), .vdd(vdd), );
  BUFX4 BUFX4_410 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf5), .Y(raddr2_0_bF_buf3_), .vdd(vdd), );
  BUFX4 BUFX4_411 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf4), .Y(raddr2_0_bF_buf2_), .vdd(vdd), );
  BUFX4 BUFX4_412 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf3), .Y(raddr2_0_bF_buf1_), .vdd(vdd), );
  BUFX4 BUFX4_413 (.gnd(gnd), .A(raddr2_0__hier0_bF_buf2), .Y(raddr2_0_bF_buf0_), .vdd(vdd), );
  BUFX4 BUFX4_414 (.gnd(gnd), .A(_2264_), .Y(_2264__bF_buf10), .vdd(vdd), );
  BUFX4 BUFX4_415 (.gnd(gnd), .A(_2264_), .Y(_2264__bF_buf9), .vdd(vdd), );
  BUFX4 BUFX4_416 (.gnd(gnd), .A(_2264_), .Y(_2264__bF_buf8), .vdd(vdd), );
  BUFX4 BUFX4_417 (.gnd(gnd), .A(_2264_), .Y(_2264__bF_buf7), .vdd(vdd), );
  BUFX4 BUFX4_418 (.gnd(gnd), .A(_2264_), .Y(_2264__bF_buf6), .vdd(vdd), );
  BUFX4 BUFX4_419 (.gnd(gnd), .A(_2264_), .Y(_2264__bF_buf5), .vdd(vdd), );
  BUFX4 BUFX4_420 (.gnd(gnd), .A(_2264_), .Y(_2264__bF_buf4), .vdd(vdd), );
  BUFX4 BUFX4_421 (.gnd(gnd), .A(_2264_), .Y(_2264__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_422 (.gnd(gnd), .A(_2264_), .Y(_2264__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_423 (.gnd(gnd), .A(_2264_), .Y(_2264__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_424 (.gnd(gnd), .A(_2264_), .Y(_2264__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_425 (.gnd(gnd), .A(_2299_), .Y(_2299__bF_buf4), .vdd(vdd), );
  BUFX4 BUFX4_426 (.gnd(gnd), .A(_2299_), .Y(_2299__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_427 (.gnd(gnd), .A(_2299_), .Y(_2299__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_428 (.gnd(gnd), .A(_2299_), .Y(_2299__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_429 (.gnd(gnd), .A(_2299_), .Y(_2299__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_430 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf96_), .vdd(vdd), );
  BUFX4 BUFX4_431 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf95_), .vdd(vdd), );
  BUFX4 BUFX4_432 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf94_), .vdd(vdd), );
  BUFX4 BUFX4_433 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf93_), .vdd(vdd), );
  BUFX4 BUFX4_434 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf92_), .vdd(vdd), );
  BUFX4 BUFX4_435 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf91_), .vdd(vdd), );
  BUFX4 BUFX4_436 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf90_), .vdd(vdd), );
  BUFX4 BUFX4_437 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf89_), .vdd(vdd), );
  BUFX4 BUFX4_438 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf88_), .vdd(vdd), );
  BUFX4 BUFX4_439 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf87_), .vdd(vdd), );
  BUFX4 BUFX4_440 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf86_), .vdd(vdd), );
  BUFX4 BUFX4_441 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf85_), .vdd(vdd), );
  BUFX4 BUFX4_442 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf84_), .vdd(vdd), );
  BUFX4 BUFX4_443 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf83_), .vdd(vdd), );
  BUFX4 BUFX4_444 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf82_), .vdd(vdd), );
  BUFX4 BUFX4_445 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf81_), .vdd(vdd), );
  BUFX4 BUFX4_446 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf80_), .vdd(vdd), );
  BUFX4 BUFX4_447 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf79_), .vdd(vdd), );
  BUFX4 BUFX4_448 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf78_), .vdd(vdd), );
  BUFX4 BUFX4_449 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf77_), .vdd(vdd), );
  BUFX4 BUFX4_450 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf76_), .vdd(vdd), );
  BUFX4 BUFX4_451 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf75_), .vdd(vdd), );
  BUFX4 BUFX4_452 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf74_), .vdd(vdd), );
  BUFX4 BUFX4_453 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf73_), .vdd(vdd), );
  BUFX4 BUFX4_454 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf72_), .vdd(vdd), );
  BUFX4 BUFX4_455 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf71_), .vdd(vdd), );
  BUFX4 BUFX4_456 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf70_), .vdd(vdd), );
  BUFX4 BUFX4_457 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf69_), .vdd(vdd), );
  BUFX4 BUFX4_458 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf68_), .vdd(vdd), );
  BUFX4 BUFX4_459 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf67_), .vdd(vdd), );
  BUFX4 BUFX4_460 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf66_), .vdd(vdd), );
  BUFX4 BUFX4_461 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf65_), .vdd(vdd), );
  BUFX4 BUFX4_462 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf64_), .vdd(vdd), );
  BUFX4 BUFX4_463 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf63_), .vdd(vdd), );
  BUFX4 BUFX4_464 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf62_), .vdd(vdd), );
  BUFX4 BUFX4_465 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf61_), .vdd(vdd), );
  BUFX4 BUFX4_466 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf60_), .vdd(vdd), );
  BUFX4 BUFX4_467 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf59_), .vdd(vdd), );
  BUFX4 BUFX4_468 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf58_), .vdd(vdd), );
  BUFX4 BUFX4_469 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf57_), .vdd(vdd), );
  BUFX4 BUFX4_470 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf56_), .vdd(vdd), );
  BUFX4 BUFX4_471 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf55_), .vdd(vdd), );
  BUFX4 BUFX4_472 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf54_), .vdd(vdd), );
  BUFX4 BUFX4_473 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf53_), .vdd(vdd), );
  BUFX4 BUFX4_474 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf52_), .vdd(vdd), );
  BUFX4 BUFX4_475 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf51_), .vdd(vdd), );
  BUFX4 BUFX4_476 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf50_), .vdd(vdd), );
  BUFX4 BUFX4_477 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf49_), .vdd(vdd), );
  BUFX4 BUFX4_478 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf48_), .vdd(vdd), );
  BUFX4 BUFX4_479 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf47_), .vdd(vdd), );
  BUFX4 BUFX4_480 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf46_), .vdd(vdd), );
  BUFX4 BUFX4_481 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf45_), .vdd(vdd), );
  BUFX4 BUFX4_482 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf44_), .vdd(vdd), );
  BUFX4 BUFX4_483 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf43_), .vdd(vdd), );
  BUFX4 BUFX4_484 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf42_), .vdd(vdd), );
  BUFX4 BUFX4_485 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf41_), .vdd(vdd), );
  BUFX4 BUFX4_486 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf40_), .vdd(vdd), );
  BUFX4 BUFX4_487 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf39_), .vdd(vdd), );
  BUFX4 BUFX4_488 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf38_), .vdd(vdd), );
  BUFX4 BUFX4_489 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf37_), .vdd(vdd), );
  BUFX4 BUFX4_490 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf36_), .vdd(vdd), );
  BUFX4 BUFX4_491 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf35_), .vdd(vdd), );
  BUFX4 BUFX4_492 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf34_), .vdd(vdd), );
  BUFX4 BUFX4_493 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf33_), .vdd(vdd), );
  BUFX4 BUFX4_494 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf32_), .vdd(vdd), );
  BUFX4 BUFX4_495 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf31_), .vdd(vdd), );
  BUFX4 BUFX4_496 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf30_), .vdd(vdd), );
  BUFX4 BUFX4_497 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf29_), .vdd(vdd), );
  BUFX4 BUFX4_498 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf28_), .vdd(vdd), );
  BUFX4 BUFX4_499 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf27_), .vdd(vdd), );
  BUFX4 BUFX4_500 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf26_), .vdd(vdd), );
  BUFX4 BUFX4_501 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf25_), .vdd(vdd), );
  BUFX4 BUFX4_502 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf24_), .vdd(vdd), );
  BUFX4 BUFX4_503 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf23_), .vdd(vdd), );
  BUFX4 BUFX4_504 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf22_), .vdd(vdd), );
  BUFX4 BUFX4_505 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf21_), .vdd(vdd), );
  BUFX4 BUFX4_506 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf20_), .vdd(vdd), );
  BUFX4 BUFX4_507 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf19_), .vdd(vdd), );
  BUFX4 BUFX4_508 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf18_), .vdd(vdd), );
  BUFX4 BUFX4_509 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf17_), .vdd(vdd), );
  BUFX4 BUFX4_510 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf16_), .vdd(vdd), );
  BUFX4 BUFX4_511 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf15_), .vdd(vdd), );
  BUFX4 BUFX4_512 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf14_), .vdd(vdd), );
  BUFX4 BUFX4_513 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf13_), .vdd(vdd), );
  BUFX4 BUFX4_514 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf12_), .vdd(vdd), );
  BUFX4 BUFX4_515 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf11_), .vdd(vdd), );
  BUFX4 BUFX4_516 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf10_), .vdd(vdd), );
  BUFX4 BUFX4_517 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf9_), .vdd(vdd), );
  BUFX4 BUFX4_518 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf8_), .vdd(vdd), );
  BUFX4 BUFX4_519 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf7_), .vdd(vdd), );
  BUFX4 BUFX4_520 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf6_), .vdd(vdd), );
  BUFX4 BUFX4_521 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf5_), .vdd(vdd), );
  BUFX4 BUFX4_522 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf4_), .vdd(vdd), );
  BUFX4 BUFX4_523 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf3_), .vdd(vdd), );
  BUFX4 BUFX4_524 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf2_), .vdd(vdd), );
  BUFX4 BUFX4_525 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf1_), .vdd(vdd), );
  BUFX4 BUFX4_526 (.gnd(gnd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf0_), .vdd(vdd), );
  BUFX4 BUFX4_527 (.gnd(gnd), .A(_1015_), .Y(_1015__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_528 (.gnd(gnd), .A(_1015_), .Y(_1015__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_529 (.gnd(gnd), .A(_1015_), .Y(_1015__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_530 (.gnd(gnd), .A(_1015_), .Y(_1015__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_531 (.gnd(gnd), .A(_1053_), .Y(_1053__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_532 (.gnd(gnd), .A(_1053_), .Y(_1053__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_533 (.gnd(gnd), .A(_1053_), .Y(_1053__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_534 (.gnd(gnd), .A(_1053_), .Y(_1053__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_535 (.gnd(gnd), .A(_992_), .Y(_992__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_536 (.gnd(gnd), .A(_992_), .Y(_992__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_537 (.gnd(gnd), .A(_992_), .Y(_992__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_538 (.gnd(gnd), .A(_992_), .Y(_992__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_539 (.gnd(gnd), .A(_2064_), .Y(_2064__bF_buf4), .vdd(vdd), );
  BUFX4 BUFX4_540 (.gnd(gnd), .A(_2064_), .Y(_2064__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_541 (.gnd(gnd), .A(_2064_), .Y(_2064__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_542 (.gnd(gnd), .A(_2064_), .Y(_2064__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_543 (.gnd(gnd), .A(_2064_), .Y(_2064__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_544 (.gnd(gnd), .A(_1009_), .Y(_1009__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_545 (.gnd(gnd), .A(_1009_), .Y(_1009__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_546 (.gnd(gnd), .A(_1009_), .Y(_1009__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_547 (.gnd(gnd), .A(_1009_), .Y(_1009__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_548 (.gnd(gnd), .A(_1047_), .Y(_1047__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_549 (.gnd(gnd), .A(_1047_), .Y(_1047__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_550 (.gnd(gnd), .A(_1047_), .Y(_1047__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_551 (.gnd(gnd), .A(_1047_), .Y(_1047__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_552 (.gnd(gnd), .A(_1141_), .Y(_1141__bF_buf7), .vdd(vdd), );
  BUFX4 BUFX4_553 (.gnd(gnd), .A(_1141_), .Y(_1141__bF_buf6), .vdd(vdd), );
  BUFX4 BUFX4_554 (.gnd(gnd), .A(_1141_), .Y(_1141__bF_buf5), .vdd(vdd), );
  BUFX4 BUFX4_555 (.gnd(gnd), .A(_1141_), .Y(_1141__bF_buf4), .vdd(vdd), );
  BUFX4 BUFX4_556 (.gnd(gnd), .A(_1141_), .Y(_1141__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_557 (.gnd(gnd), .A(_1141_), .Y(_1141__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_558 (.gnd(gnd), .A(_1141_), .Y(_1141__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_559 (.gnd(gnd), .A(_1141_), .Y(_1141__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_560 (.gnd(gnd), .A(_1902_), .Y(_1902__bF_buf7), .vdd(vdd), );
  BUFX4 BUFX4_561 (.gnd(gnd), .A(_1902_), .Y(_1902__bF_buf6), .vdd(vdd), );
  BUFX4 BUFX4_562 (.gnd(gnd), .A(_1902_), .Y(_1902__bF_buf5), .vdd(vdd), );
  BUFX4 BUFX4_563 (.gnd(gnd), .A(_1902_), .Y(_1902__bF_buf4), .vdd(vdd), );
  BUFX4 BUFX4_564 (.gnd(gnd), .A(_1902_), .Y(_1902__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_565 (.gnd(gnd), .A(_1902_), .Y(_1902__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_566 (.gnd(gnd), .A(_1902_), .Y(_1902__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_567 (.gnd(gnd), .A(_1902_), .Y(_1902__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_568 (.gnd(gnd), .A(_1003_), .Y(_1003__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_569 (.gnd(gnd), .A(_1003_), .Y(_1003__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_570 (.gnd(gnd), .A(_1003_), .Y(_1003__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_571 (.gnd(gnd), .A(_1003_), .Y(_1003__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_572 (.gnd(gnd), .A(_1041_), .Y(_1041__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_573 (.gnd(gnd), .A(_1041_), .Y(_1041__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_574 (.gnd(gnd), .A(_1041_), .Y(_1041__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_575 (.gnd(gnd), .A(_1041_), .Y(_1041__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_576 (.gnd(gnd), .A(_1000_), .Y(_1000__bF_buf7), .vdd(vdd), );
  BUFX4 BUFX4_577 (.gnd(gnd), .A(_1000_), .Y(_1000__bF_buf6), .vdd(vdd), );
  BUFX4 BUFX4_578 (.gnd(gnd), .A(_1000_), .Y(_1000__bF_buf5), .vdd(vdd), );
  BUFX4 BUFX4_579 (.gnd(gnd), .A(_1000_), .Y(_1000__bF_buf4), .vdd(vdd), );
  BUFX4 BUFX4_580 (.gnd(gnd), .A(_1000_), .Y(_1000__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_581 (.gnd(gnd), .A(_1000_), .Y(_1000__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_582 (.gnd(gnd), .A(_1000_), .Y(_1000__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_583 (.gnd(gnd), .A(_1000_), .Y(_1000__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_584 (.gnd(gnd), .A(_1705_), .Y(_1705__bF_buf7), .vdd(vdd), );
  BUFX4 BUFX4_585 (.gnd(gnd), .A(_1705_), .Y(_1705__bF_buf6), .vdd(vdd), );
  BUFX4 BUFX4_586 (.gnd(gnd), .A(_1705_), .Y(_1705__bF_buf5), .vdd(vdd), );
  BUFX4 BUFX4_587 (.gnd(gnd), .A(_1705_), .Y(_1705__bF_buf4), .vdd(vdd), );
  BUFX4 BUFX4_588 (.gnd(gnd), .A(_1705_), .Y(_1705__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_589 (.gnd(gnd), .A(_1705_), .Y(_1705__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_590 (.gnd(gnd), .A(_1705_), .Y(_1705__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_591 (.gnd(gnd), .A(_1705_), .Y(_1705__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_592 (.gnd(gnd), .A(_1035_), .Y(_1035__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_593 (.gnd(gnd), .A(_1035_), .Y(_1035__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_594 (.gnd(gnd), .A(_1035_), .Y(_1035__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_595 (.gnd(gnd), .A(_1035_), .Y(_1035__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_596 (.gnd(gnd), .A(_1605_), .Y(_1605__bF_buf7), .vdd(vdd), );
  BUFX4 BUFX4_597 (.gnd(gnd), .A(_1605_), .Y(_1605__bF_buf6), .vdd(vdd), );
  BUFX4 BUFX4_598 (.gnd(gnd), .A(_1605_), .Y(_1605__bF_buf5), .vdd(vdd), );
  BUFX4 BUFX4_599 (.gnd(gnd), .A(_1605_), .Y(_1605__bF_buf4), .vdd(vdd), );
  BUFX4 BUFX4_600 (.gnd(gnd), .A(_1605_), .Y(_1605__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_601 (.gnd(gnd), .A(_1605_), .Y(_1605__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_602 (.gnd(gnd), .A(_1605_), .Y(_1605__bF_buf1), .vdd(vdd), );
  BUFX4 BUFX4_603 (.gnd(gnd), .A(_1605_), .Y(_1605__bF_buf0), .vdd(vdd), );
  BUFX4 BUFX4_604 (.gnd(gnd), .A(_1070_), .Y(_1070__bF_buf10), .vdd(vdd), );
  BUFX4 BUFX4_605 (.gnd(gnd), .A(_1070_), .Y(_1070__bF_buf9), .vdd(vdd), );
  BUFX4 BUFX4_606 (.gnd(gnd), .A(_1070_), .Y(_1070__bF_buf8), .vdd(vdd), );
  BUFX4 BUFX4_607 (.gnd(gnd), .A(_1070_), .Y(_1070__bF_buf7), .vdd(vdd), );
  BUFX4 BUFX4_608 (.gnd(gnd), .A(_1070_), .Y(_1070__bF_buf6), .vdd(vdd), );
  BUFX4 BUFX4_609 (.gnd(gnd), .A(_1070_), .Y(_1070__bF_buf5), .vdd(vdd), );
  BUFX4 BUFX4_610 (.gnd(gnd), .A(_1070_), .Y(_1070__bF_buf4), .vdd(vdd), );
  BUFX4 BUFX4_611 (.gnd(gnd), .A(_1070_), .Y(_1070__bF_buf3), .vdd(vdd), );
  BUFX4 BUFX4_612 (.gnd(gnd), .A(_1070_), .Y(_1070__bF_buf2), .vdd(vdd), );
  BUFX4 BUFX4_613 (.Y(_1070__bF_buf1), .A(_1070_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_614 (.Y(_1070__bF_buf0), .A(_1070_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_615 (.Y(_1966__bF_buf7), .A(_1966_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_616 (.Y(_1966__bF_buf6), .A(_1966_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_617 (.Y(_1966__bF_buf5), .A(_1966_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_618 (.Y(_1966__bF_buf4), .A(_1966_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_619 (.Y(_1966__bF_buf3), .A(_1966_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_620 (.Y(_1966__bF_buf2), .A(_1966_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_621 (.Y(_1966__bF_buf1), .A(_1966_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_622 (.Y(_1966__bF_buf0), .A(_1966_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_623 (.Y(_1029__bF_buf3), .A(_1029_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_624 (.Y(_1029__bF_buf2), .A(_1029_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_625 (.Y(_1029__bF_buf1), .A(_1029_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_626 (.Y(_1029__bF_buf0), .A(_1029_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_627 (.Y(_4036__bF_buf8), .A(_4036_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_628 (.Y(_4036__bF_buf7), .A(_4036_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_629 (.Y(_4036__bF_buf6), .A(_4036_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_630 (.Y(_4036__bF_buf5), .A(_4036_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_631 (.Y(_4036__bF_buf4), .A(_4036_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_632 (.Y(_4036__bF_buf3), .A(_4036_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_633 (.Y(_4036__bF_buf2), .A(_4036_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_634 (.Y(_4036__bF_buf1), .A(_4036_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_635 (.Y(_4036__bF_buf0), .A(_4036_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_636 (.Y(_1408__bF_buf7), .A(_1408_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_637 (.Y(_1408__bF_buf6), .A(_1408_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_638 (.Y(_1408__bF_buf5), .A(_1408_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_639 (.Y(_1408__bF_buf4), .A(_1408_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_640 (.Y(_1408__bF_buf3), .A(_1408_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_641 (.Y(_1408__bF_buf2), .A(_1408_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_642 (.Y(_1408__bF_buf1), .A(_1408_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_643 (.Y(_1408__bF_buf0), .A(_1408_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_644 (.Y(_1769__bF_buf7), .A(_1769_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_645 (.Y(_1769__bF_buf6), .A(_1769_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_646 (.Y(_1769__bF_buf5), .A(_1769_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_647 (.Y(_1769__bF_buf4), .A(_1769_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_648 (.Y(_1769__bF_buf3), .A(_1769_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_649 (.Y(_1769__bF_buf2), .A(_1769_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_650 (.Y(_1769__bF_buf1), .A(_1769_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_651 (.Y(_1769__bF_buf0), .A(_1769_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_652 (.Y(_4033__bF_buf7), .A(_4033_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_653 (.Y(_4033__bF_buf6), .A(_4033_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_654 (.Y(_4033__bF_buf5), .A(_4033_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_655 (.Y(_4033__bF_buf4), .A(_4033_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_656 (.Y(_4033__bF_buf3), .A(_4033_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_657 (.Y(_4033__bF_buf2), .A(_4033_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_658 (.Y(_4033__bF_buf1), .A(_4033_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_659 (.Y(_4033__bF_buf0), .A(_4033_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_660 (.Y(_2231__bF_buf4), .A(_2231_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_661 (.Y(_2231__bF_buf3), .A(_2231_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_662 (.Y(_2231__bF_buf2), .A(_2231_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_663 (.Y(_2231__bF_buf1), .A(_2231_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_664 (.Y(_2231__bF_buf0), .A(_2231_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_665 (.Y(_1023__bF_buf3), .A(_1023_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_666 (.Y(_1023__bF_buf2), .A(_1023_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_667 (.Y(_1023__bF_buf1), .A(_1023_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_668 (.Y(_1023__bF_buf0), .A(_1023_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_669 (.Y(raddr2_2_bF_buf10_), .A(raddr2[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_670 (.Y(raddr2_2_bF_buf9_), .A(raddr2[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_671 (.Y(raddr2_2_bF_buf8_), .A(raddr2[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_672 (.Y(raddr2_2_bF_buf7_), .A(raddr2[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_673 (.Y(raddr2_2_bF_buf6_), .A(raddr2[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_674 (.Y(raddr2_2_bF_buf5_), .A(raddr2[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_675 (.Y(raddr2_2_bF_buf4_), .A(raddr2[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_676 (.Y(raddr2_2_bF_buf3_), .A(raddr2[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_677 (.Y(raddr2_2_bF_buf2_), .A(raddr2[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_678 (.Y(raddr2_2_bF_buf1_), .A(raddr2[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_679 (.Y(raddr2_2_bF_buf0_), .A(raddr2[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_680 (.Y(_1061__bF_buf3), .A(_1061_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_681 (.Y(_1061__bF_buf2), .A(_1061_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_682 (.Y(_1061__bF_buf1), .A(_1061_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_683 (.Y(_1061__bF_buf0), .A(_1061_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_684 (.Y(_2398__bF_buf7), .A(_2398_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_685 (.Y(_2398__bF_buf6), .A(_2398_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_686 (.Y(_2398__bF_buf5), .A(_2398_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_687 (.Y(_2398__bF_buf4), .A(_2398_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_688 (.Y(_2398__bF_buf3), .A(_2398_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_689 (.Y(_2398__bF_buf2), .A(_2398_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_690 (.Y(_2398__bF_buf1), .A(_2398_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_691 (.Y(_2398__bF_buf0), .A(_2398_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_692 (.Y(_1669__bF_buf4), .A(_1669_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_693 (.Y(_1669__bF_buf3), .A(_1669_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_694 (.Y(_1669__bF_buf2), .A(_1669_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_695 (.Y(_1669__bF_buf1), .A(_1669_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_696 (.Y(_1669__bF_buf0), .A(_1669_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_697 (.Y(raddr1_2_bF_buf10_), .A(raddr1[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_698 (.Y(raddr1_2_bF_buf9_), .A(raddr1[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_699 (.Y(raddr1_2_bF_buf8_), .A(raddr1[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_700 (.Y(raddr1_2_bF_buf7_), .A(raddr1[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_701 (.Y(raddr1_2_bF_buf6_), .A(raddr1[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_702 (.Y(raddr1_2_bF_buf5_), .A(raddr1[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_703 (.Y(raddr1_2_bF_buf4_), .A(raddr1[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_704 (.Y(raddr1_2_bF_buf3_), .A(raddr1[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_705 (.Y(raddr1_2_bF_buf2_), .A(raddr1[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_706 (.Y(raddr1_2_bF_buf1_), .A(raddr1[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_707 (.Y(raddr1_2_bF_buf0_), .A(raddr1[2]), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_708 (.Y(_1017__bF_buf3), .A(_1017_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_709 (.Y(_1017__bF_buf2), .A(_1017_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_710 (.Y(_1017__bF_buf1), .A(_1017_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_711 (.Y(_1017__bF_buf0), .A(_1017_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_712 (.Y(_1055__bF_buf3), .A(_1055_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_713 (.Y(_1055__bF_buf2), .A(_1055_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_714 (.Y(_1055__bF_buf1), .A(_1055_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_715 (.Y(_1055__bF_buf0), .A(_1055_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_716 (.Y(_1472__bF_buf4), .A(_1472_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_717 (.Y(_1472__bF_buf3), .A(_1472_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_718 (.Y(_1472__bF_buf2), .A(_1472_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_719 (.Y(_1472__bF_buf1), .A(_1472_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_720 (.Y(_1472__bF_buf0), .A(_1472_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_721 (.Y(_2198__bF_buf4), .A(_2198_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_722 (.Y(_2198__bF_buf3), .A(_2198_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_723 (.Y(_2198__bF_buf2), .A(_2198_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_724 (.Y(_2198__bF_buf1), .A(_2198_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_725 (.Y(_2198__bF_buf0), .A(_2198_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_726 (.Y(_1049__bF_buf3), .A(_1049_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_727 (.Y(_1049__bF_buf2), .A(_1049_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_728 (.Y(_1049__bF_buf1), .A(_1049_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_729 (.Y(_1049__bF_buf0), .A(_1049_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_730 (.Y(_1011__bF_buf3), .A(_1011_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_731 (.Y(_1011__bF_buf2), .A(_1011_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_732 (.Y(_1011__bF_buf1), .A(_1011_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_733 (.Y(_1011__bF_buf0), .A(_1011_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_734 (.Y(_1240__bF_buf4), .A(_1240_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_735 (.Y(_1240__bF_buf3), .A(_1240_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_736 (.Y(_1240__bF_buf2), .A(_1240_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_737 (.Y(_1240__bF_buf1), .A(_1240_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_738 (.Y(_1240__bF_buf0), .A(_1240_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_739 (.Y(_1105__bF_buf7), .A(_1105_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_740 (.Y(_1105__bF_buf6), .A(_1105_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_741 (.Y(_1105__bF_buf5), .A(_1105_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_742 (.Y(_1105__bF_buf4), .A(_1105_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_743 (.Y(_1105__bF_buf3), .A(_1105_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_744 (.Y(_1105__bF_buf2), .A(_1105_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_745 (.Y(_1105__bF_buf1), .A(_1105_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_746 (.Y(_1105__bF_buf0), .A(_1105_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_747 (.Y(_1143__bF_buf7), .A(_1143_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_748 (.Y(_1143__bF_buf6), .A(_1143_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_749 (.Y(_1143__bF_buf5), .A(_1143_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_750 (.Y(_1143__bF_buf4), .A(_1143_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_751 (.Y(_1143__bF_buf3), .A(_1143_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_752 (.Y(_1143__bF_buf2), .A(_1143_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_753 (.Y(_1143__bF_buf1), .A(_1143_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_754 (.Y(_1143__bF_buf0), .A(_1143_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_755 (.Y(_1005__bF_buf3), .A(_1005_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_756 (.Y(_1005__bF_buf2), .A(_1005_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_757 (.Y(_1005__bF_buf1), .A(_1005_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_758 (.Y(_1005__bF_buf0), .A(_1005_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_759 (.Y(_1043__bF_buf3), .A(_1043_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_760 (.Y(_1043__bF_buf2), .A(_1043_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_761 (.Y(_1043__bF_buf1), .A(_1043_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_762 (.Y(_1043__bF_buf0), .A(_1043_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_763 (.Y(_1901__bF_buf5), .A(_1901_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_764 (.Y(_1901__bF_buf4), .A(_1901_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_765 (.Y(_1901__bF_buf3), .A(_1901_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_766 (.Y(_1901__bF_buf2), .A(_1901_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_767 (.Y(_1901__bF_buf1), .A(_1901_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_768 (.Y(_1901__bF_buf0), .A(_1901_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_769 (.Y(_1037__bF_buf3), .A(_1037_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_770 (.Y(_1037__bF_buf2), .A(_1037_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_771 (.Y(_1037__bF_buf1), .A(_1037_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_772 (.Y(_1037__bF_buf0), .A(_1037_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_773 (.Y(_1704__bF_buf5), .A(_1704_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_774 (.Y(_1704__bF_buf4), .A(_1704_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_775 (.Y(_1704__bF_buf3), .A(_1704_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_776 (.Y(_1704__bF_buf2), .A(_1704_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_777 (.Y(_1704__bF_buf1), .A(_1704_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_778 (.Y(_1704__bF_buf0), .A(_1704_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_779 (.Y(_1069__bF_buf4), .A(_1069_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_780 (.Y(_1069__bF_buf3), .A(_1069_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_781 (.Y(_1069__bF_buf2), .A(_1069_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_782 (.Y(_1069__bF_buf1), .A(_1069_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_783 (.Y(_1069__bF_buf0), .A(_1069_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_784 (.Y(_4038__bF_buf8), .A(_4038_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_785 (.Y(_4038__bF_buf7), .A(_4038_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_786 (.Y(_4038__bF_buf6), .A(_4038_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_787 (.Y(_4038__bF_buf5), .A(_4038_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_788 (.Y(_4038__bF_buf4), .A(_4038_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_789 (.Y(_4038__bF_buf3), .A(_4038_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_790 (.Y(_4038__bF_buf2), .A(_4038_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_791 (.Y(_4038__bF_buf1), .A(_4038_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_792 (.Y(_4038__bF_buf0), .A(_4038_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_793 (.Y(_1031__bF_buf3), .A(_1031_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_794 (.Y(_1031__bF_buf2), .A(_1031_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_795 (.Y(_1031__bF_buf1), .A(_1031_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_796 (.Y(_1031__bF_buf0), .A(_1031_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_797 (.Y(_1507__bF_buf7), .A(_1507_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_798 (.Y(_1507__bF_buf6), .A(_1507_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_799 (.Y(_1507__bF_buf5), .A(_1507_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_800 (.Y(_1507__bF_buf4), .A(_1507_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_801 (.Y(_1507__bF_buf3), .A(_1507_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_802 (.Y(_1507__bF_buf2), .A(_1507_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_803 (.Y(_1507__bF_buf1), .A(_1507_), .gnd(gnd), .vdd(vdd), );
  BUFX4 BUFX4_804 (.Y(_1507__bF_buf0), .A(_1507_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1 (.Y(_1279_), .A(_1141__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf14), .C(regs_24__4_), );
  OAI21X1 OAI21X1_2 (.Y(_538_), .A(_1274__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1009__bF_buf3), .C(_1279_), );
  OAI21X1 OAI21X1_3 (.Y(_1280_), .A(_1141__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf13), .C(regs_24__5_), );
  OAI21X1 OAI21X1_4 (.Y(_539_), .A(_1274__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1011__bF_buf3), .C(_1280_), );
  OAI21X1 OAI21X1_5 (.Y(_1281_), .A(_1141__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf12), .C(regs_24__6_), );
  OAI21X1 OAI21X1_6 (.Y(_540_), .A(_1274__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1013__bF_buf3), .C(_1281_), );
  OAI21X1 OAI21X1_7 (.Y(_1282_), .A(_1141__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf11), .C(regs_24__7_), );
  OAI21X1 OAI21X1_8 (.Y(_541_), .A(_1274__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1015__bF_buf3), .C(_1282_), );
  OAI21X1 OAI21X1_9 (.Y(_1283_), .A(_1141__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf10), .C(regs_24__8_), );
  OAI21X1 OAI21X1_10 (.Y(_542_), .A(_1274__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1017__bF_buf3), .C(_1283_), );
  OAI21X1 OAI21X1_11 (.Y(_1284_), .A(_1141__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf9), .C(regs_24__9_), );
  OAI21X1 OAI21X1_12 (.Y(_543_), .A(_1274__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1019__bF_buf3), .C(_1284_), );
  OAI21X1 OAI21X1_13 (.Y(_1285_), .A(_1141__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf8), .C(regs_24__10_), );
  OAI21X1 OAI21X1_14 (.Y(_513_), .A(_1274__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1021__bF_buf3), .C(_1285_), );
  OAI21X1 OAI21X1_15 (.Y(_1286_), .A(_1141__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf7), .C(regs_24__11_), );
  OAI21X1 OAI21X1_16 (.Y(_514_), .A(_1274__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1023__bF_buf3), .C(_1286_), );
  OAI21X1 OAI21X1_17 (.Y(_1287_), .A(_1141__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf6), .C(regs_24__12_), );
  OAI21X1 OAI21X1_18 (.Y(_515_), .A(_1274__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1025__bF_buf3), .C(_1287_), );
  OAI21X1 OAI21X1_19 (.Y(_1288_), .A(_1141__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf5), .C(regs_24__13_), );
  OAI21X1 OAI21X1_20 (.Y(_516_), .A(_1274__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1027__bF_buf3), .C(_1288_), );
  OAI21X1 OAI21X1_21 (.Y(_1289_), .A(_1141__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf4), .C(regs_24__14_), );
  OAI21X1 OAI21X1_22 (.Y(_517_), .A(_1274__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1029__bF_buf3), .C(_1289_), );
  OAI21X1 OAI21X1_23 (.Y(_1290_), .A(_1141__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf3), .C(regs_24__15_), );
  OAI21X1 OAI21X1_24 (.Y(_518_), .A(_1274__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1031__bF_buf3), .C(_1290_), );
  OAI21X1 OAI21X1_25 (.Y(_1291_), .A(_1141__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf2), .C(regs_24__16_), );
  OAI21X1 OAI21X1_26 (.Y(_519_), .A(_1274__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1033__bF_buf3), .C(_1291_), );
  OAI21X1 OAI21X1_27 (.Y(_1292_), .A(_1141__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf1), .C(regs_24__17_), );
  OAI21X1 OAI21X1_28 (.Y(_520_), .A(_1274__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1035__bF_buf3), .C(_1292_), );
  OAI21X1 OAI21X1_29 (.Y(_1293_), .A(_1141__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf0), .C(regs_24__18_), );
  OAI21X1 OAI21X1_30 (.Y(_521_), .A(_1274__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1037__bF_buf3), .C(_1293_), );
  OAI21X1 OAI21X1_31 (.Y(_1294_), .A(_1141__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf14), .C(regs_24__19_), );
  OAI21X1 OAI21X1_32 (.Y(_522_), .A(_1274__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1039__bF_buf3), .C(_1294_), );
  OAI21X1 OAI21X1_33 (.Y(_1295_), .A(_1141__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf13), .C(regs_24__20_), );
  OAI21X1 OAI21X1_34 (.Y(_524_), .A(_1274__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1041__bF_buf3), .C(_1295_), );
  OAI21X1 OAI21X1_35 (.Y(_1296_), .A(_1141__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf12), .C(regs_24__21_), );
  OAI21X1 OAI21X1_36 (.Y(_525_), .A(_1274__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1043__bF_buf3), .C(_1296_), );
  OAI21X1 OAI21X1_37 (.Y(_1297_), .A(_1141__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf11), .C(regs_24__22_), );
  OAI21X1 OAI21X1_38 (.Y(_526_), .A(_1274__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1045__bF_buf3), .C(_1297_), );
  OAI21X1 OAI21X1_39 (.Y(_1298_), .A(_1141__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf10), .C(regs_24__23_), );
  OAI21X1 OAI21X1_40 (.Y(_527_), .A(_1274__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1047__bF_buf3), .C(_1298_), );
  OAI21X1 OAI21X1_41 (.Y(_1299_), .A(_1141__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf9), .C(regs_24__24_), );
  OAI21X1 OAI21X1_42 (.Y(_528_), .A(_1274__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1049__bF_buf3), .C(_1299_), );
  OAI21X1 OAI21X1_43 (.Y(_1300_), .A(_1141__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf8), .C(regs_24__25_), );
  OAI21X1 OAI21X1_44 (.Y(_529_), .A(_1274__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1051__bF_buf3), .C(_1300_), );
  OAI21X1 OAI21X1_45 (.Y(_1301_), .A(_1141__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf7), .C(regs_24__26_), );
  OAI21X1 OAI21X1_46 (.Y(_530_), .A(_1274__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1053__bF_buf3), .C(_1301_), );
  OAI21X1 OAI21X1_47 (.Y(_1302_), .A(_1141__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf6), .C(regs_24__27_), );
  OAI21X1 OAI21X1_48 (.Y(_531_), .A(_1274__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1055__bF_buf3), .C(_1302_), );
  OAI21X1 OAI21X1_49 (.Y(_1303_), .A(_1141__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf5), .C(regs_24__28_), );
  OAI21X1 OAI21X1_50 (.Y(_532_), .A(_1274__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1057__bF_buf3), .C(_1303_), );
  OAI21X1 OAI21X1_51 (.Y(_1304_), .A(_1141__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf4), .C(regs_24__29_), );
  OAI21X1 OAI21X1_52 (.Y(_533_), .A(_1274__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1059__bF_buf3), .C(_1304_), );
  OAI21X1 OAI21X1_53 (.Y(_1305_), .A(_1141__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf3), .C(regs_24__30_), );
  OAI21X1 OAI21X1_54 (.Y(_535_), .A(_1274__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1061__bF_buf3), .C(_1305_), );
  OAI21X1 OAI21X1_55 (.Y(_1306_), .A(_1141__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf2), .C(regs_24__31_), );
  OAI21X1 OAI21X1_56 (.Y(_536_), .A(_1274__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1063__bF_buf3), .C(_1306_), );
  INVX2 INVX2_1 (.Y(_1307_), .A(regs_23__0_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_1 (.Y(_1308_), .A(waddr[3]), .gnd(gnd), .vdd(vdd), .B(_993_), );
  OR2X2 OR2X2_1 (.Y(_1309_), .A(_1308_), .gnd(gnd), .vdd(vdd), .B(waddr[2]), );
  NOR2X1 NOR2X1_1 (.Y(_1310_), .A(_1142__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_1309__bF_buf5), );
  NAND2X1 NAND2X1_2 (.Y(_1311_), .A(wdata[0]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf7), );
  OAI21X1 OAI21X1_57 (.Y(_480_), .A(_1307_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf6), .C(_1311_), );
  INVX2 INVX2_2 (.Y(_1312_), .A(regs_23__1_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_3 (.Y(_1313_), .A(wdata[1]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf5), );
  OAI21X1 OAI21X1_58 (.Y(_491_), .A(_1312_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf4), .C(_1313_), );
  INVX2 INVX2_3 (.Y(_1314_), .A(regs_23__2_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_4 (.Y(_1315_), .A(wdata[2]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf3), );
  OAI21X1 OAI21X1_59 (.Y(_502_), .A(_1314_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf2), .C(_1315_), );
  INVX2 INVX2_4 (.Y(_1316_), .A(regs_23__3_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_5 (.Y(_1317_), .A(wdata[3]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf1), );
  OAI21X1 OAI21X1_60 (.Y(_505_), .A(_1316_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf0), .C(_1317_), );
  INVX2 INVX2_5 (.Y(_1318_), .A(regs_23__4_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_6 (.Y(_1319_), .A(wdata[4]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf7), );
  OAI21X1 OAI21X1_61 (.Y(_506_), .A(_1318_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf6), .C(_1319_), );
  INVX2 INVX2_6 (.Y(_1320_), .A(regs_23__5_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_7 (.Y(_1321_), .A(wdata[5]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf5), );
  OAI21X1 OAI21X1_62 (.Y(_507_), .A(_1320_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf4), .C(_1321_), );
  INVX2 INVX2_7 (.Y(_1322_), .A(regs_23__6_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_8 (.Y(_1323_), .A(wdata[6]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf3), );
  OAI21X1 OAI21X1_63 (.Y(_508_), .A(_1322_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf2), .C(_1323_), );
  INVX2 INVX2_8 (.Y(_1324_), .A(regs_23__7_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_9 (.Y(_1325_), .A(wdata[7]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf1), );
  OAI21X1 OAI21X1_64 (.Y(_509_), .A(_1324_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf0), .C(_1325_), );
  INVX2 INVX2_9 (.Y(_1326_), .A(regs_23__8_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_10 (.Y(_1327_), .A(wdata[8]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf7), );
  OAI21X1 OAI21X1_65 (.Y(_510_), .A(_1326_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf6), .C(_1327_), );
  INVX2 INVX2_10 (.Y(_1328_), .A(regs_23__9_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_11 (.Y(_1329_), .A(wdata[9]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf5), );
  OAI21X1 OAI21X1_66 (.Y(_511_), .A(_1328_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf4), .C(_1329_), );
  INVX2 INVX2_11 (.Y(_1330_), .A(regs_23__10_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_12 (.Y(_1331_), .A(wdata[10]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf3), );
  OAI21X1 OAI21X1_67 (.Y(_481_), .A(_1330_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf2), .C(_1331_), );
  INVX2 INVX2_12 (.Y(_1332_), .A(regs_23__11_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_13 (.Y(_1333_), .A(wdata[11]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf1), );
  OAI21X1 OAI21X1_68 (.Y(_482_), .A(_1332_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf0), .C(_1333_), );
  INVX2 INVX2_13 (.Y(_1334_), .A(regs_23__12_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_14 (.Y(_1335_), .A(wdata[12]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf7), );
  OAI21X1 OAI21X1_69 (.Y(_483_), .A(_1334_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf6), .C(_1335_), );
  INVX2 INVX2_14 (.Y(_1336_), .A(regs_23__13_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_15 (.Y(_1337_), .A(wdata[13]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf5), );
  OAI21X1 OAI21X1_70 (.Y(_484_), .A(_1336_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf4), .C(_1337_), );
  INVX2 INVX2_15 (.Y(_1338_), .A(regs_23__14_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_16 (.Y(_1339_), .A(wdata[14]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf3), );
  OAI21X1 OAI21X1_71 (.Y(_485_), .A(_1338_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf2), .C(_1339_), );
  INVX2 INVX2_16 (.Y(_1340_), .A(regs_23__15_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_17 (.Y(_1341_), .A(wdata[15]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf1), );
  OAI21X1 OAI21X1_72 (.Y(_486_), .A(_1340_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf0), .C(_1341_), );
  INVX2 INVX2_17 (.Y(_1342_), .A(regs_23__16_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_18 (.Y(_1343_), .A(wdata[16]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf7), );
  OAI21X1 OAI21X1_73 (.Y(_487_), .A(_1342_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf6), .C(_1343_), );
  INVX2 INVX2_18 (.Y(_1344_), .A(regs_23__17_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_19 (.Y(_1345_), .A(wdata[17]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf5), );
  OAI21X1 OAI21X1_74 (.Y(_488_), .A(_1344_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf4), .C(_1345_), );
  INVX2 INVX2_19 (.Y(_1346_), .A(regs_23__18_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_20 (.Y(_1347_), .A(wdata[18]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf3), );
  OAI21X1 OAI21X1_75 (.Y(_489_), .A(_1346_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf2), .C(_1347_), );
  INVX2 INVX2_20 (.Y(_1348_), .A(regs_23__19_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_21 (.Y(_1349_), .A(wdata[19]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf1), );
  OAI21X1 OAI21X1_76 (.Y(_490_), .A(_1348_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf0), .C(_1349_), );
  INVX2 INVX2_21 (.Y(_1350_), .A(regs_23__20_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_22 (.Y(_1351_), .A(wdata[20]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf7), );
  OAI21X1 OAI21X1_77 (.Y(_492_), .A(_1350_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf6), .C(_1351_), );
  INVX2 INVX2_22 (.Y(_1352_), .A(regs_23__21_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_23 (.Y(_1353_), .A(wdata[21]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf5), );
  OAI21X1 OAI21X1_78 (.Y(_493_), .A(_1352_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf4), .C(_1353_), );
  INVX2 INVX2_23 (.Y(_1354_), .A(regs_23__22_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_24 (.Y(_1355_), .A(wdata[22]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf3), );
  OAI21X1 OAI21X1_79 (.Y(_494_), .A(_1354_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf2), .C(_1355_), );
  INVX2 INVX2_24 (.Y(_1356_), .A(regs_23__23_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_25 (.Y(_1357_), .A(wdata[23]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf1), );
  OAI21X1 OAI21X1_80 (.Y(_495_), .A(_1356_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf0), .C(_1357_), );
  INVX2 INVX2_25 (.Y(_1358_), .A(regs_23__24_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_26 (.Y(_1359_), .A(wdata[24]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf7), );
  OAI21X1 OAI21X1_81 (.Y(_496_), .A(_1358_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf6), .C(_1359_), );
  INVX2 INVX2_26 (.Y(_1360_), .A(regs_23__25_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_27 (.Y(_1361_), .A(wdata[25]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf5), );
  OAI21X1 OAI21X1_82 (.Y(_497_), .A(_1360_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf4), .C(_1361_), );
  INVX2 INVX2_27 (.Y(_1362_), .A(regs_23__26_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_28 (.Y(_1363_), .A(wdata[26]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf3), );
  OAI21X1 OAI21X1_83 (.Y(_498_), .A(_1362_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf2), .C(_1363_), );
  INVX2 INVX2_28 (.Y(_1364_), .A(regs_23__27_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_29 (.Y(_1365_), .A(wdata[27]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf1), );
  OAI21X1 OAI21X1_84 (.Y(_499_), .A(_1364_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf0), .C(_1365_), );
  INVX2 INVX2_29 (.Y(_1366_), .A(regs_23__28_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_30 (.Y(_1367_), .A(wdata[28]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf7), );
  OAI21X1 OAI21X1_85 (.Y(_500_), .A(_1366_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf6), .C(_1367_), );
  INVX2 INVX2_30 (.Y(_1368_), .A(regs_23__29_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_31 (.Y(_1369_), .A(wdata[29]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf5), );
  OAI21X1 OAI21X1_86 (.Y(_501_), .A(_1368_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf4), .C(_1369_), );
  INVX2 INVX2_31 (.Y(_1370_), .A(regs_23__30_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_32 (.Y(_1371_), .A(wdata[30]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf3), );
  OAI21X1 OAI21X1_87 (.Y(_503_), .A(_1370_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf2), .C(_1371_), );
  INVX2 INVX2_32 (.Y(_1372_), .A(regs_23__31_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_33 (.Y(_1373_), .A(wdata[31]), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf1), );
  OAI21X1 OAI21X1_88 (.Y(_504_), .A(_1372_), .gnd(gnd), .vdd(vdd), .B(_1310__bF_buf0), .C(_1373_), );
  NOR2X1 NOR2X1_2 (.Y(_1374_), .A(_1001__bF_buf9), .gnd(gnd), .vdd(vdd), .B(_1309__bF_buf4), );
  NOR2X1 NOR2X1_3 (.Y(_1375_), .A(regs_22__0_), .gnd(gnd), .vdd(vdd), .B(_1374__bF_buf7), );
  AOI21X1 AOI21X1_1 (.Y(_448_), .A(_992__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1374__bF_buf6), .C(_1375_), );
  NOR2X1 NOR2X1_4 (.Y(_1376_), .A(regs_22__1_), .gnd(gnd), .vdd(vdd), .B(_1374__bF_buf5), );
  AOI21X1 AOI21X1_2 (.Y(_459_), .A(_1003__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1374__bF_buf4), .C(_1376_), );
  NOR2X1 NOR2X1_5 (.Y(_1377_), .A(regs_22__2_), .gnd(gnd), .vdd(vdd), .B(_1374__bF_buf3), );
  AOI21X1 AOI21X1_3 (.Y(_470_), .A(_1005__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1374__bF_buf2), .C(_1377_), );
  NOR2X1 NOR2X1_6 (.Y(_1378_), .A(regs_22__3_), .gnd(gnd), .vdd(vdd), .B(_1374__bF_buf1), );
  AOI21X1 AOI21X1_4 (.gnd(gnd), .A(_1007__bF_buf3), .Y(_473_), .vdd(vdd), .B(_1374__bF_buf0), .C(_1378_), );
  NOR2X1 NOR2X1_7 (.gnd(gnd), .A(regs_22__4_), .Y(_1379_), .vdd(vdd), .B(_1374__bF_buf7), );
  AOI21X1 AOI21X1_5 (.gnd(gnd), .A(_1009__bF_buf2), .Y(_474_), .vdd(vdd), .B(_1374__bF_buf6), .C(_1379_), );
  NOR2X1 NOR2X1_8 (.gnd(gnd), .A(regs_22__5_), .Y(_1380_), .vdd(vdd), .B(_1374__bF_buf5), );
  AOI21X1 AOI21X1_6 (.gnd(gnd), .A(_1011__bF_buf2), .Y(_475_), .vdd(vdd), .B(_1374__bF_buf4), .C(_1380_), );
  NOR2X1 NOR2X1_9 (.gnd(gnd), .A(regs_22__6_), .Y(_1381_), .vdd(vdd), .B(_1374__bF_buf3), );
  AOI21X1 AOI21X1_7 (.gnd(gnd), .A(_1013__bF_buf2), .Y(_476_), .vdd(vdd), .B(_1374__bF_buf2), .C(_1381_), );
  NOR2X1 NOR2X1_10 (.gnd(gnd), .A(regs_22__7_), .Y(_1382_), .vdd(vdd), .B(_1374__bF_buf1), );
  AOI21X1 AOI21X1_8 (.gnd(gnd), .A(_1015__bF_buf2), .Y(_477_), .vdd(vdd), .B(_1374__bF_buf0), .C(_1382_), );
  NOR2X1 NOR2X1_11 (.gnd(gnd), .A(regs_22__8_), .Y(_1383_), .vdd(vdd), .B(_1374__bF_buf7), );
  AOI21X1 AOI21X1_9 (.gnd(gnd), .A(_1017__bF_buf2), .Y(_478_), .vdd(vdd), .B(_1374__bF_buf6), .C(_1383_), );
  NOR2X1 NOR2X1_12 (.gnd(gnd), .A(regs_22__9_), .Y(_1384_), .vdd(vdd), .B(_1374__bF_buf5), );
  AOI21X1 AOI21X1_10 (.gnd(gnd), .A(_1019__bF_buf2), .Y(_479_), .vdd(vdd), .B(_1374__bF_buf4), .C(_1384_), );
  NOR2X1 NOR2X1_13 (.gnd(gnd), .A(regs_22__10_), .Y(_1385_), .vdd(vdd), .B(_1374__bF_buf3), );
  AOI21X1 AOI21X1_11 (.gnd(gnd), .A(_1021__bF_buf2), .Y(_449_), .vdd(vdd), .B(_1374__bF_buf2), .C(_1385_), );
  NOR2X1 NOR2X1_14 (.gnd(gnd), .A(regs_22__11_), .Y(_1386_), .vdd(vdd), .B(_1374__bF_buf1), );
  AOI21X1 AOI21X1_12 (.gnd(gnd), .A(_1023__bF_buf2), .Y(_450_), .vdd(vdd), .B(_1374__bF_buf0), .C(_1386_), );
  NOR2X1 NOR2X1_15 (.gnd(gnd), .A(regs_22__12_), .Y(_1387_), .vdd(vdd), .B(_1374__bF_buf7), );
  AOI21X1 AOI21X1_13 (.gnd(gnd), .A(_1025__bF_buf2), .Y(_451_), .vdd(vdd), .B(_1374__bF_buf6), .C(_1387_), );
  NOR2X1 NOR2X1_16 (.gnd(gnd), .A(regs_22__13_), .Y(_1388_), .vdd(vdd), .B(_1374__bF_buf5), );
  AOI21X1 AOI21X1_14 (.gnd(gnd), .A(_1027__bF_buf2), .Y(_452_), .vdd(vdd), .B(_1374__bF_buf4), .C(_1388_), );
  NOR2X1 NOR2X1_17 (.gnd(gnd), .A(regs_22__14_), .Y(_1389_), .vdd(vdd), .B(_1374__bF_buf3), );
  AOI21X1 AOI21X1_15 (.gnd(gnd), .A(_1029__bF_buf2), .Y(_453_), .vdd(vdd), .B(_1374__bF_buf2), .C(_1389_), );
  NOR2X1 NOR2X1_18 (.gnd(gnd), .A(regs_22__15_), .Y(_1390_), .vdd(vdd), .B(_1374__bF_buf1), );
  AOI21X1 AOI21X1_16 (.gnd(gnd), .A(_1031__bF_buf2), .Y(_454_), .vdd(vdd), .B(_1374__bF_buf0), .C(_1390_), );
  NOR2X1 NOR2X1_19 (.gnd(gnd), .A(regs_22__16_), .Y(_1391_), .vdd(vdd), .B(_1374__bF_buf7), );
  AOI21X1 AOI21X1_17 (.gnd(gnd), .A(_1033__bF_buf2), .Y(_455_), .vdd(vdd), .B(_1374__bF_buf6), .C(_1391_), );
  NOR2X1 NOR2X1_20 (.gnd(gnd), .A(regs_22__17_), .Y(_1392_), .vdd(vdd), .B(_1374__bF_buf5), );
  AOI21X1 AOI21X1_18 (.gnd(gnd), .A(_1035__bF_buf2), .Y(_456_), .vdd(vdd), .B(_1374__bF_buf4), .C(_1392_), );
  NOR2X1 NOR2X1_21 (.gnd(gnd), .A(regs_22__18_), .Y(_1393_), .vdd(vdd), .B(_1374__bF_buf3), );
  AOI21X1 AOI21X1_19 (.gnd(gnd), .A(_1037__bF_buf2), .Y(_457_), .vdd(vdd), .B(_1374__bF_buf2), .C(_1393_), );
  NOR2X1 NOR2X1_22 (.gnd(gnd), .A(regs_22__19_), .Y(_1394_), .vdd(vdd), .B(_1374__bF_buf1), );
  AOI21X1 AOI21X1_20 (.gnd(gnd), .A(_1039__bF_buf2), .Y(_458_), .vdd(vdd), .B(_1374__bF_buf0), .C(_1394_), );
  NOR2X1 NOR2X1_23 (.gnd(gnd), .A(regs_22__20_), .Y(_1395_), .vdd(vdd), .B(_1374__bF_buf7), );
  AOI21X1 AOI21X1_21 (.gnd(gnd), .A(_1041__bF_buf2), .Y(_460_), .vdd(vdd), .B(_1374__bF_buf6), .C(_1395_), );
  NOR2X1 NOR2X1_24 (.gnd(gnd), .A(regs_22__21_), .Y(_1396_), .vdd(vdd), .B(_1374__bF_buf5), );
  AOI21X1 AOI21X1_22 (.gnd(gnd), .A(_1043__bF_buf2), .Y(_461_), .vdd(vdd), .B(_1374__bF_buf4), .C(_1396_), );
  NOR2X1 NOR2X1_25 (.gnd(gnd), .A(regs_22__22_), .Y(_1397_), .vdd(vdd), .B(_1374__bF_buf3), );
  AOI21X1 AOI21X1_23 (.gnd(gnd), .A(_1045__bF_buf2), .Y(_462_), .vdd(vdd), .B(_1374__bF_buf2), .C(_1397_), );
  NOR2X1 NOR2X1_26 (.gnd(gnd), .A(regs_22__23_), .Y(_1398_), .vdd(vdd), .B(_1374__bF_buf1), );
  AOI21X1 AOI21X1_24 (.gnd(gnd), .A(_1047__bF_buf2), .Y(_463_), .vdd(vdd), .B(_1374__bF_buf0), .C(_1398_), );
  NOR2X1 NOR2X1_27 (.gnd(gnd), .A(regs_22__24_), .Y(_1399_), .vdd(vdd), .B(_1374__bF_buf7), );
  AOI21X1 AOI21X1_25 (.gnd(gnd), .A(_1049__bF_buf2), .Y(_464_), .vdd(vdd), .B(_1374__bF_buf6), .C(_1399_), );
  NOR2X1 NOR2X1_28 (.gnd(gnd), .A(regs_22__25_), .Y(_1400_), .vdd(vdd), .B(_1374__bF_buf5), );
  AOI21X1 AOI21X1_26 (.gnd(gnd), .A(_1051__bF_buf2), .Y(_465_), .vdd(vdd), .B(_1374__bF_buf4), .C(_1400_), );
  NOR2X1 NOR2X1_29 (.gnd(gnd), .A(regs_22__26_), .Y(_1401_), .vdd(vdd), .B(_1374__bF_buf3), );
  AOI21X1 AOI21X1_27 (.gnd(gnd), .A(_1053__bF_buf2), .Y(_466_), .vdd(vdd), .B(_1374__bF_buf2), .C(_1401_), );
  NOR2X1 NOR2X1_30 (.gnd(gnd), .A(regs_22__27_), .Y(_1402_), .vdd(vdd), .B(_1374__bF_buf1), );
  AOI21X1 AOI21X1_28 (.gnd(gnd), .A(_1055__bF_buf2), .Y(_467_), .vdd(vdd), .B(_1374__bF_buf0), .C(_1402_), );
  NOR2X1 NOR2X1_31 (.gnd(gnd), .A(regs_22__28_), .Y(_1403_), .vdd(vdd), .B(_1374__bF_buf7), );
  AOI21X1 AOI21X1_29 (.gnd(gnd), .A(_1057__bF_buf2), .Y(_468_), .vdd(vdd), .B(_1374__bF_buf6), .C(_1403_), );
  NOR2X1 NOR2X1_32 (.gnd(gnd), .A(regs_22__29_), .Y(_1404_), .vdd(vdd), .B(_1374__bF_buf5), );
  AOI21X1 AOI21X1_30 (.gnd(gnd), .A(_1059__bF_buf2), .Y(_469_), .vdd(vdd), .B(_1374__bF_buf4), .C(_1404_), );
  NOR2X1 NOR2X1_33 (.gnd(gnd), .A(regs_22__30_), .Y(_1405_), .vdd(vdd), .B(_1374__bF_buf3), );
  AOI21X1 AOI21X1_31 (.gnd(gnd), .A(_1061__bF_buf2), .Y(_471_), .vdd(vdd), .B(_1374__bF_buf2), .C(_1405_), );
  NOR2X1 NOR2X1_34 (.gnd(gnd), .A(regs_22__31_), .Y(_1406_), .vdd(vdd), .B(_1374__bF_buf1), );
  AOI21X1 AOI21X1_32 (.gnd(gnd), .A(_1063__bF_buf2), .Y(_472_), .vdd(vdd), .B(_1374__bF_buf0), .C(_1406_), );
  INVX2 INVX2_33 (.gnd(gnd), .A(regs_21__0_), .Y(_1407_), .vdd(vdd), );
  NOR2X1 NOR2X1_35 (.gnd(gnd), .A(_1309__bF_buf3), .Y(_1408_), .vdd(vdd), .B(_1070__bF_buf10), );
  NAND2X1 NAND2X1_34 (.gnd(gnd), .A(wdata[0]), .Y(_1409_), .vdd(vdd), .B(_1408__bF_buf7), );
  OAI21X1 OAI21X1_89 (.gnd(gnd), .A(_1407_), .Y(_416_), .vdd(vdd), .B(_1408__bF_buf6), .C(_1409_), );
  INVX2 INVX2_34 (.gnd(gnd), .A(regs_21__1_), .Y(_1410_), .vdd(vdd), );
  NAND2X1 NAND2X1_35 (.gnd(gnd), .A(wdata[1]), .Y(_1411_), .vdd(vdd), .B(_1408__bF_buf5), );
  OAI21X1 OAI21X1_90 (.gnd(gnd), .A(_1410_), .Y(_427_), .vdd(vdd), .B(_1408__bF_buf4), .C(_1411_), );
  INVX2 INVX2_35 (.gnd(gnd), .A(regs_21__2_), .Y(_1412_), .vdd(vdd), );
  NAND2X1 NAND2X1_36 (.gnd(gnd), .A(wdata[2]), .Y(_1413_), .vdd(vdd), .B(_1408__bF_buf3), );
  OAI21X1 OAI21X1_91 (.gnd(gnd), .A(_1412_), .Y(_438_), .vdd(vdd), .B(_1408__bF_buf2), .C(_1413_), );
  INVX2 INVX2_36 (.gnd(gnd), .A(regs_21__3_), .Y(_1414_), .vdd(vdd), );
  NAND2X1 NAND2X1_37 (.gnd(gnd), .A(wdata[3]), .Y(_1415_), .vdd(vdd), .B(_1408__bF_buf1), );
  OAI21X1 OAI21X1_92 (.gnd(gnd), .A(_1414_), .Y(_441_), .vdd(vdd), .B(_1408__bF_buf0), .C(_1415_), );
  INVX2 INVX2_37 (.gnd(gnd), .A(regs_21__4_), .Y(_1416_), .vdd(vdd), );
  NAND2X1 NAND2X1_38 (.gnd(gnd), .A(wdata[4]), .Y(_1417_), .vdd(vdd), .B(_1408__bF_buf7), );
  OAI21X1 OAI21X1_93 (.gnd(gnd), .A(_1416_), .Y(_442_), .vdd(vdd), .B(_1408__bF_buf6), .C(_1417_), );
  INVX2 INVX2_38 (.gnd(gnd), .A(regs_21__5_), .Y(_1418_), .vdd(vdd), );
  NAND2X1 NAND2X1_39 (.gnd(gnd), .A(wdata[5]), .Y(_1419_), .vdd(vdd), .B(_1408__bF_buf5), );
  OAI21X1 OAI21X1_94 (.gnd(gnd), .A(_1418_), .Y(_443_), .vdd(vdd), .B(_1408__bF_buf4), .C(_1419_), );
  INVX2 INVX2_39 (.gnd(gnd), .A(regs_21__6_), .Y(_1420_), .vdd(vdd), );
  NAND2X1 NAND2X1_40 (.gnd(gnd), .A(wdata[6]), .Y(_1421_), .vdd(vdd), .B(_1408__bF_buf3), );
  OAI21X1 OAI21X1_95 (.gnd(gnd), .A(_1420_), .Y(_444_), .vdd(vdd), .B(_1408__bF_buf2), .C(_1421_), );
  INVX2 INVX2_40 (.gnd(gnd), .A(regs_21__7_), .Y(_1422_), .vdd(vdd), );
  NAND2X1 NAND2X1_41 (.gnd(gnd), .A(wdata[7]), .Y(_1423_), .vdd(vdd), .B(_1408__bF_buf1), );
  OAI21X1 OAI21X1_96 (.gnd(gnd), .A(_1422_), .Y(_445_), .vdd(vdd), .B(_1408__bF_buf0), .C(_1423_), );
  INVX2 INVX2_41 (.gnd(gnd), .A(regs_21__8_), .Y(_1424_), .vdd(vdd), );
  NAND2X1 NAND2X1_42 (.gnd(gnd), .A(wdata[8]), .Y(_1425_), .vdd(vdd), .B(_1408__bF_buf7), );
  OAI21X1 OAI21X1_97 (.gnd(gnd), .A(_1424_), .Y(_446_), .vdd(vdd), .B(_1408__bF_buf6), .C(_1425_), );
  INVX2 INVX2_42 (.gnd(gnd), .A(regs_21__9_), .Y(_1426_), .vdd(vdd), );
  NAND2X1 NAND2X1_43 (.gnd(gnd), .A(wdata[9]), .Y(_1427_), .vdd(vdd), .B(_1408__bF_buf5), );
  OAI21X1 OAI21X1_98 (.gnd(gnd), .A(_1426_), .Y(_447_), .vdd(vdd), .B(_1408__bF_buf4), .C(_1427_), );
  INVX2 INVX2_43 (.gnd(gnd), .A(regs_21__10_), .Y(_1428_), .vdd(vdd), );
  NAND2X1 NAND2X1_44 (.gnd(gnd), .A(wdata[10]), .Y(_1429_), .vdd(vdd), .B(_1408__bF_buf3), );
  OAI21X1 OAI21X1_99 (.gnd(gnd), .A(_1428_), .Y(_417_), .vdd(vdd), .B(_1408__bF_buf2), .C(_1429_), );
  INVX2 INVX2_44 (.gnd(gnd), .A(regs_21__11_), .Y(_1430_), .vdd(vdd), );
  NAND2X1 NAND2X1_45 (.gnd(gnd), .A(wdata[11]), .Y(_1431_), .vdd(vdd), .B(_1408__bF_buf1), );
  OAI21X1 OAI21X1_100 (.gnd(gnd), .A(_1430_), .Y(_418_), .vdd(vdd), .B(_1408__bF_buf0), .C(_1431_), );
  INVX2 INVX2_45 (.gnd(gnd), .A(regs_21__12_), .Y(_1432_), .vdd(vdd), );
  NAND2X1 NAND2X1_46 (.gnd(gnd), .A(wdata[12]), .Y(_1433_), .vdd(vdd), .B(_1408__bF_buf7), );
  OAI21X1 OAI21X1_101 (.gnd(gnd), .A(_1432_), .Y(_419_), .vdd(vdd), .B(_1408__bF_buf6), .C(_1433_), );
  INVX2 INVX2_46 (.gnd(gnd), .A(regs_21__13_), .Y(_1434_), .vdd(vdd), );
  NAND2X1 NAND2X1_47 (.gnd(gnd), .A(wdata[13]), .Y(_1435_), .vdd(vdd), .B(_1408__bF_buf5), );
  OAI21X1 OAI21X1_102 (.gnd(gnd), .A(_1434_), .Y(_420_), .vdd(vdd), .B(_1408__bF_buf4), .C(_1435_), );
  INVX2 INVX2_47 (.gnd(gnd), .A(regs_21__14_), .Y(_1436_), .vdd(vdd), );
  NAND2X1 NAND2X1_48 (.gnd(gnd), .A(wdata[14]), .Y(_1437_), .vdd(vdd), .B(_1408__bF_buf3), );
  OAI21X1 OAI21X1_103 (.gnd(gnd), .A(_1436_), .Y(_421_), .vdd(vdd), .B(_1408__bF_buf2), .C(_1437_), );
  INVX2 INVX2_48 (.gnd(gnd), .A(regs_21__15_), .Y(_1438_), .vdd(vdd), );
  NAND2X1 NAND2X1_49 (.gnd(gnd), .A(wdata[15]), .Y(_1439_), .vdd(vdd), .B(_1408__bF_buf1), );
  OAI21X1 OAI21X1_104 (.gnd(gnd), .A(_1438_), .Y(_422_), .vdd(vdd), .B(_1408__bF_buf0), .C(_1439_), );
  INVX2 INVX2_49 (.gnd(gnd), .A(regs_21__16_), .Y(_1440_), .vdd(vdd), );
  NAND2X1 NAND2X1_50 (.gnd(gnd), .A(wdata[16]), .Y(_1441_), .vdd(vdd), .B(_1408__bF_buf7), );
  OAI21X1 OAI21X1_105 (.gnd(gnd), .A(_1440_), .Y(_423_), .vdd(vdd), .B(_1408__bF_buf6), .C(_1441_), );
  INVX2 INVX2_50 (.gnd(gnd), .A(regs_21__17_), .Y(_1442_), .vdd(vdd), );
  NAND2X1 NAND2X1_51 (.gnd(gnd), .A(wdata[17]), .Y(_1443_), .vdd(vdd), .B(_1408__bF_buf5), );
  OAI21X1 OAI21X1_106 (.gnd(gnd), .A(_1442_), .Y(_424_), .vdd(vdd), .B(_1408__bF_buf4), .C(_1443_), );
  INVX2 INVX2_51 (.gnd(gnd), .A(regs_21__18_), .Y(_1444_), .vdd(vdd), );
  NAND2X1 NAND2X1_52 (.gnd(gnd), .A(wdata[18]), .Y(_1445_), .vdd(vdd), .B(_1408__bF_buf3), );
  OAI21X1 OAI21X1_107 (.gnd(gnd), .A(_1444_), .Y(_425_), .vdd(vdd), .B(_1408__bF_buf2), .C(_1445_), );
  INVX2 INVX2_52 (.gnd(gnd), .A(regs_21__19_), .Y(_1446_), .vdd(vdd), );
  NAND2X1 NAND2X1_53 (.gnd(gnd), .A(wdata[19]), .Y(_1447_), .vdd(vdd), .B(_1408__bF_buf1), );
  OAI21X1 OAI21X1_108 (.gnd(gnd), .A(_1446_), .Y(_426_), .vdd(vdd), .B(_1408__bF_buf0), .C(_1447_), );
  INVX2 INVX2_53 (.gnd(gnd), .A(regs_21__20_), .Y(_1448_), .vdd(vdd), );
  NAND2X1 NAND2X1_54 (.gnd(gnd), .A(wdata[20]), .Y(_1449_), .vdd(vdd), .B(_1408__bF_buf7), );
  OAI21X1 OAI21X1_109 (.gnd(gnd), .A(_1448_), .Y(_428_), .vdd(vdd), .B(_1408__bF_buf6), .C(_1449_), );
  INVX2 INVX2_54 (.gnd(gnd), .A(regs_21__21_), .Y(_1450_), .vdd(vdd), );
  NAND2X1 NAND2X1_55 (.gnd(gnd), .A(wdata[21]), .Y(_1451_), .vdd(vdd), .B(_1408__bF_buf5), );
  OAI21X1 OAI21X1_110 (.gnd(gnd), .A(_1450_), .Y(_429_), .vdd(vdd), .B(_1408__bF_buf4), .C(_1451_), );
  INVX2 INVX2_55 (.gnd(gnd), .A(regs_21__22_), .Y(_1452_), .vdd(vdd), );
  NAND2X1 NAND2X1_56 (.gnd(gnd), .A(wdata[22]), .Y(_1453_), .vdd(vdd), .B(_1408__bF_buf3), );
  OAI21X1 OAI21X1_111 (.gnd(gnd), .A(_1452_), .Y(_430_), .vdd(vdd), .B(_1408__bF_buf2), .C(_1453_), );
  INVX2 INVX2_56 (.gnd(gnd), .A(regs_21__23_), .Y(_1454_), .vdd(vdd), );
  NAND2X1 NAND2X1_57 (.gnd(gnd), .A(wdata[23]), .Y(_1455_), .vdd(vdd), .B(_1408__bF_buf1), );
  OAI21X1 OAI21X1_112 (.gnd(gnd), .A(_1454_), .Y(_431_), .vdd(vdd), .B(_1408__bF_buf0), .C(_1455_), );
  INVX2 INVX2_57 (.gnd(gnd), .A(regs_21__24_), .Y(_1456_), .vdd(vdd), );
  NAND2X1 NAND2X1_58 (.gnd(gnd), .A(wdata[24]), .Y(_1457_), .vdd(vdd), .B(_1408__bF_buf7), );
  OAI21X1 OAI21X1_113 (.gnd(gnd), .A(_1456_), .Y(_432_), .vdd(vdd), .B(_1408__bF_buf6), .C(_1457_), );
  INVX2 INVX2_58 (.gnd(gnd), .A(regs_21__25_), .Y(_1458_), .vdd(vdd), );
  NAND2X1 NAND2X1_59 (.gnd(gnd), .A(wdata[25]), .Y(_1459_), .vdd(vdd), .B(_1408__bF_buf5), );
  OAI21X1 OAI21X1_114 (.gnd(gnd), .A(_1458_), .Y(_433_), .vdd(vdd), .B(_1408__bF_buf4), .C(_1459_), );
  INVX2 INVX2_59 (.gnd(gnd), .A(regs_21__26_), .Y(_1460_), .vdd(vdd), );
  NAND2X1 NAND2X1_60 (.gnd(gnd), .A(wdata[26]), .Y(_1461_), .vdd(vdd), .B(_1408__bF_buf3), );
  OAI21X1 OAI21X1_115 (.gnd(gnd), .A(_1460_), .Y(_434_), .vdd(vdd), .B(_1408__bF_buf2), .C(_1461_), );
  INVX2 INVX2_60 (.gnd(gnd), .A(regs_21__27_), .Y(_1462_), .vdd(vdd), );
  NAND2X1 NAND2X1_61 (.gnd(gnd), .A(wdata[27]), .Y(_1463_), .vdd(vdd), .B(_1408__bF_buf1), );
  OAI21X1 OAI21X1_116 (.gnd(gnd), .A(_1462_), .Y(_435_), .vdd(vdd), .B(_1408__bF_buf0), .C(_1463_), );
  INVX2 INVX2_61 (.gnd(gnd), .A(regs_21__28_), .Y(_1464_), .vdd(vdd), );
  NAND2X1 NAND2X1_62 (.gnd(gnd), .A(wdata[28]), .Y(_1465_), .vdd(vdd), .B(_1408__bF_buf7), );
  OAI21X1 OAI21X1_117 (.gnd(gnd), .A(_1464_), .Y(_436_), .vdd(vdd), .B(_1408__bF_buf6), .C(_1465_), );
  INVX2 INVX2_62 (.gnd(gnd), .A(regs_21__29_), .Y(_1466_), .vdd(vdd), );
  NAND2X1 NAND2X1_63 (.gnd(gnd), .A(wdata[29]), .Y(_1467_), .vdd(vdd), .B(_1408__bF_buf5), );
  OAI21X1 OAI21X1_118 (.gnd(gnd), .A(_1466_), .Y(_437_), .vdd(vdd), .B(_1408__bF_buf4), .C(_1467_), );
  INVX2 INVX2_63 (.gnd(gnd), .A(regs_21__30_), .Y(_1468_), .vdd(vdd), );
  NAND2X1 NAND2X1_64 (.gnd(gnd), .A(wdata[30]), .Y(_1469_), .vdd(vdd), .B(_1408__bF_buf3), );
  OAI21X1 OAI21X1_119 (.gnd(gnd), .A(_1468_), .Y(_439_), .vdd(vdd), .B(_1408__bF_buf2), .C(_1469_), );
  INVX2 INVX2_64 (.gnd(gnd), .A(regs_21__31_), .Y(_1470_), .vdd(vdd), );
  NAND2X1 NAND2X1_65 (.gnd(gnd), .A(wdata[31]), .Y(_1471_), .vdd(vdd), .B(_1408__bF_buf1), );
  OAI21X1 OAI21X1_120 (.gnd(gnd), .A(_1470_), .Y(_440_), .vdd(vdd), .B(_1408__bF_buf0), .C(_1471_), );
  OR2X2 OR2X2_2 (.gnd(gnd), .A(_1309__bF_buf2), .Y(_1472_), .vdd(vdd), .B(_1104__bF_buf1), );
  OAI21X1 OAI21X1_121 (.gnd(gnd), .A(_1309__bF_buf1), .Y(_1473_), .vdd(vdd), .B(_1104__bF_buf0), .C(regs_20__0_), );
  OAI21X1 OAI21X1_122 (.gnd(gnd), .A(_1472__bF_buf4), .Y(_384_), .vdd(vdd), .B(_992__bF_buf2), .C(_1473_), );
  OAI21X1 OAI21X1_123 (.gnd(gnd), .A(_1309__bF_buf0), .Y(_1474_), .vdd(vdd), .B(_1104__bF_buf14), .C(regs_20__1_), );
  OAI21X1 OAI21X1_124 (.gnd(gnd), .A(_1472__bF_buf3), .Y(_395_), .vdd(vdd), .B(_1003__bF_buf2), .C(_1474_), );
  OAI21X1 OAI21X1_125 (.gnd(gnd), .A(_1309__bF_buf5), .Y(_1475_), .vdd(vdd), .B(_1104__bF_buf13), .C(regs_20__2_), );
  OAI21X1 OAI21X1_126 (.gnd(gnd), .A(_1472__bF_buf2), .Y(_406_), .vdd(vdd), .B(_1005__bF_buf2), .C(_1475_), );
  OAI21X1 OAI21X1_127 (.gnd(gnd), .A(_1309__bF_buf4), .Y(_1476_), .vdd(vdd), .B(_1104__bF_buf12), .C(regs_20__3_), );
  OAI21X1 OAI21X1_128 (.gnd(gnd), .A(_1472__bF_buf1), .Y(_409_), .vdd(vdd), .B(_1007__bF_buf2), .C(_1476_), );
  OAI21X1 OAI21X1_129 (.gnd(gnd), .A(_1309__bF_buf3), .Y(_1477_), .vdd(vdd), .B(_1104__bF_buf11), .C(regs_20__4_), );
  OAI21X1 OAI21X1_130 (.gnd(gnd), .A(_1472__bF_buf0), .Y(_410_), .vdd(vdd), .B(_1009__bF_buf1), .C(_1477_), );
  OAI21X1 OAI21X1_131 (.gnd(gnd), .A(_1309__bF_buf2), .Y(_1478_), .vdd(vdd), .B(_1104__bF_buf10), .C(regs_20__5_), );
  OAI21X1 OAI21X1_132 (.gnd(gnd), .A(_1472__bF_buf4), .Y(_411_), .vdd(vdd), .B(_1011__bF_buf1), .C(_1478_), );
  OAI21X1 OAI21X1_133 (.gnd(gnd), .A(_1309__bF_buf1), .Y(_1479_), .vdd(vdd), .B(_1104__bF_buf9), .C(regs_20__6_), );
  OAI21X1 OAI21X1_134 (.gnd(gnd), .A(_1472__bF_buf3), .Y(_412_), .vdd(vdd), .B(_1013__bF_buf1), .C(_1479_), );
  OAI21X1 OAI21X1_135 (.gnd(gnd), .A(_1309__bF_buf0), .Y(_1480_), .vdd(vdd), .B(_1104__bF_buf8), .C(regs_20__7_), );
  OAI21X1 OAI21X1_136 (.gnd(gnd), .A(_1472__bF_buf2), .Y(_413_), .vdd(vdd), .B(_1015__bF_buf1), .C(_1480_), );
  OAI21X1 OAI21X1_137 (.gnd(gnd), .A(_1309__bF_buf5), .Y(_1481_), .vdd(vdd), .B(_1104__bF_buf7), .C(regs_20__8_), );
  OAI21X1 OAI21X1_138 (.gnd(gnd), .A(_1472__bF_buf1), .Y(_414_), .vdd(vdd), .B(_1017__bF_buf1), .C(_1481_), );
  OAI21X1 OAI21X1_139 (.gnd(gnd), .A(_1309__bF_buf4), .Y(_1482_), .vdd(vdd), .B(_1104__bF_buf6), .C(regs_20__9_), );
  OAI21X1 OAI21X1_140 (.gnd(gnd), .A(_1472__bF_buf0), .Y(_415_), .vdd(vdd), .B(_1019__bF_buf1), .C(_1482_), );
  OAI21X1 OAI21X1_141 (.gnd(gnd), .A(_1309__bF_buf3), .Y(_1483_), .vdd(vdd), .B(_1104__bF_buf5), .C(regs_20__10_), );
  OAI21X1 OAI21X1_142 (.gnd(gnd), .A(_1472__bF_buf4), .Y(_385_), .vdd(vdd), .B(_1021__bF_buf1), .C(_1483_), );
  OAI21X1 OAI21X1_143 (.gnd(gnd), .A(_1309__bF_buf2), .Y(_1484_), .vdd(vdd), .B(_1104__bF_buf4), .C(regs_20__11_), );
  OAI21X1 OAI21X1_144 (.gnd(gnd), .A(_1472__bF_buf3), .Y(_386_), .vdd(vdd), .B(_1023__bF_buf1), .C(_1484_), );
  OAI21X1 OAI21X1_145 (.gnd(gnd), .A(_1309__bF_buf1), .Y(_1485_), .vdd(vdd), .B(_1104__bF_buf3), .C(regs_20__12_), );
  OAI21X1 OAI21X1_146 (.gnd(gnd), .A(_1472__bF_buf2), .Y(_387_), .vdd(vdd), .B(_1025__bF_buf1), .C(_1485_), );
  OAI21X1 OAI21X1_147 (.gnd(gnd), .A(_1309__bF_buf0), .Y(_1486_), .vdd(vdd), .B(_1104__bF_buf2), .C(regs_20__13_), );
  OAI21X1 OAI21X1_148 (.gnd(gnd), .A(_1472__bF_buf1), .Y(_388_), .vdd(vdd), .B(_1027__bF_buf1), .C(_1486_), );
  OAI21X1 OAI21X1_149 (.gnd(gnd), .A(_1309__bF_buf5), .Y(_1487_), .vdd(vdd), .B(_1104__bF_buf1), .C(regs_20__14_), );
  OAI21X1 OAI21X1_150 (.gnd(gnd), .A(_1472__bF_buf0), .Y(_389_), .vdd(vdd), .B(_1029__bF_buf1), .C(_1487_), );
  OAI21X1 OAI21X1_151 (.gnd(gnd), .A(_1309__bF_buf4), .Y(_1488_), .vdd(vdd), .B(_1104__bF_buf0), .C(regs_20__15_), );
  OAI21X1 OAI21X1_152 (.gnd(gnd), .A(_1472__bF_buf4), .Y(_390_), .vdd(vdd), .B(_1031__bF_buf1), .C(_1488_), );
  OAI21X1 OAI21X1_153 (.gnd(gnd), .A(_1309__bF_buf3), .Y(_1489_), .vdd(vdd), .B(_1104__bF_buf14), .C(regs_20__16_), );
  OAI21X1 OAI21X1_154 (.gnd(gnd), .A(_1472__bF_buf3), .Y(_391_), .vdd(vdd), .B(_1033__bF_buf1), .C(_1489_), );
  OAI21X1 OAI21X1_155 (.gnd(gnd), .A(_1309__bF_buf2), .Y(_1490_), .vdd(vdd), .B(_1104__bF_buf13), .C(regs_20__17_), );
  OAI21X1 OAI21X1_156 (.gnd(gnd), .A(_1472__bF_buf2), .Y(_392_), .vdd(vdd), .B(_1035__bF_buf1), .C(_1490_), );
  OAI21X1 OAI21X1_157 (.gnd(gnd), .A(_1309__bF_buf1), .Y(_1491_), .vdd(vdd), .B(_1104__bF_buf12), .C(regs_20__18_), );
  OAI21X1 OAI21X1_158 (.gnd(gnd), .A(_1472__bF_buf1), .Y(_393_), .vdd(vdd), .B(_1037__bF_buf1), .C(_1491_), );
  OAI21X1 OAI21X1_159 (.gnd(gnd), .A(_1309__bF_buf0), .Y(_1492_), .vdd(vdd), .B(_1104__bF_buf11), .C(regs_20__19_), );
  OAI21X1 OAI21X1_160 (.gnd(gnd), .A(_1472__bF_buf0), .Y(_394_), .vdd(vdd), .B(_1039__bF_buf1), .C(_1492_), );
  OAI21X1 OAI21X1_161 (.gnd(gnd), .A(_1309__bF_buf5), .Y(_1493_), .vdd(vdd), .B(_1104__bF_buf10), .C(regs_20__20_), );
  OAI21X1 OAI21X1_162 (.gnd(gnd), .A(_1472__bF_buf4), .Y(_396_), .vdd(vdd), .B(_1041__bF_buf1), .C(_1493_), );
  OAI21X1 OAI21X1_163 (.gnd(gnd), .A(_1309__bF_buf4), .Y(_1494_), .vdd(vdd), .B(_1104__bF_buf9), .C(regs_20__21_), );
  OAI21X1 OAI21X1_164 (.gnd(gnd), .A(_1472__bF_buf3), .Y(_397_), .vdd(vdd), .B(_1043__bF_buf1), .C(_1494_), );
  OAI21X1 OAI21X1_165 (.gnd(gnd), .A(_1309__bF_buf3), .Y(_1495_), .vdd(vdd), .B(_1104__bF_buf8), .C(regs_20__22_), );
  OAI21X1 OAI21X1_166 (.gnd(gnd), .A(_1472__bF_buf2), .Y(_398_), .vdd(vdd), .B(_1045__bF_buf1), .C(_1495_), );
  OAI21X1 OAI21X1_167 (.gnd(gnd), .A(_1309__bF_buf2), .Y(_1496_), .vdd(vdd), .B(_1104__bF_buf7), .C(regs_20__23_), );
  OAI21X1 OAI21X1_168 (.gnd(gnd), .A(_1472__bF_buf1), .Y(_399_), .vdd(vdd), .B(_1047__bF_buf1), .C(_1496_), );
  OAI21X1 OAI21X1_169 (.gnd(gnd), .A(_1309__bF_buf1), .Y(_1497_), .vdd(vdd), .B(_1104__bF_buf6), .C(regs_20__24_), );
  OAI21X1 OAI21X1_170 (.gnd(gnd), .A(_1472__bF_buf0), .Y(_400_), .vdd(vdd), .B(_1049__bF_buf1), .C(_1497_), );
  OAI21X1 OAI21X1_171 (.gnd(gnd), .A(_1309__bF_buf0), .Y(_1498_), .vdd(vdd), .B(_1104__bF_buf5), .C(regs_20__25_), );
  OAI21X1 OAI21X1_172 (.gnd(gnd), .A(_1472__bF_buf4), .Y(_401_), .vdd(vdd), .B(_1051__bF_buf1), .C(_1498_), );
  OAI21X1 OAI21X1_173 (.gnd(gnd), .A(_1309__bF_buf5), .Y(_1499_), .vdd(vdd), .B(_1104__bF_buf4), .C(regs_20__26_), );
  OAI21X1 OAI21X1_174 (.gnd(gnd), .A(_1472__bF_buf3), .Y(_402_), .vdd(vdd), .B(_1053__bF_buf1), .C(_1499_), );
  OAI21X1 OAI21X1_175 (.gnd(gnd), .A(_1309__bF_buf4), .Y(_1500_), .vdd(vdd), .B(_1104__bF_buf3), .C(regs_20__27_), );
  OAI21X1 OAI21X1_176 (.gnd(gnd), .A(_1472__bF_buf2), .Y(_403_), .vdd(vdd), .B(_1055__bF_buf1), .C(_1500_), );
  OAI21X1 OAI21X1_177 (.gnd(gnd), .A(_1309__bF_buf3), .Y(_1501_), .vdd(vdd), .B(_1104__bF_buf2), .C(regs_20__28_), );
  OAI21X1 OAI21X1_178 (.gnd(gnd), .A(_1472__bF_buf1), .Y(_404_), .vdd(vdd), .B(_1057__bF_buf1), .C(_1501_), );
  OAI21X1 OAI21X1_179 (.gnd(gnd), .A(_1309__bF_buf2), .Y(_1502_), .vdd(vdd), .B(_1104__bF_buf1), .C(regs_20__29_), );
  OAI21X1 OAI21X1_180 (.gnd(gnd), .A(_1472__bF_buf0), .Y(_405_), .vdd(vdd), .B(_1059__bF_buf1), .C(_1502_), );
  OAI21X1 OAI21X1_181 (.gnd(gnd), .A(_1309__bF_buf1), .Y(_1503_), .vdd(vdd), .B(_1104__bF_buf0), .C(regs_20__30_), );
  OAI21X1 OAI21X1_182 (.gnd(gnd), .A(_1472__bF_buf4), .Y(_407_), .vdd(vdd), .B(_1061__bF_buf1), .C(_1503_), );
  OAI21X1 OAI21X1_183 (.gnd(gnd), .A(_1309__bF_buf0), .Y(_1504_), .vdd(vdd), .B(_1104__bF_buf14), .C(regs_20__31_), );
  OAI21X1 OAI21X1_184 (.gnd(gnd), .A(_1472__bF_buf3), .Y(_408_), .vdd(vdd), .B(_1063__bF_buf1), .C(_1504_), );
  INVX2 INVX2_65 (.gnd(gnd), .A(regs_19__0_), .Y(_1505_), .vdd(vdd), );
  OR2X2 OR2X2_3 (.gnd(gnd), .A(_1308_), .Y(_1506_), .vdd(vdd), .B(_1139_), );
  NOR2X1 NOR2X1_36 (.gnd(gnd), .A(_1142__bF_buf4), .Y(_1507_), .vdd(vdd), .B(_1506__bF_buf5), );
  NAND2X1 NAND2X1_66 (.gnd(gnd), .A(wdata[0]), .Y(_1508_), .vdd(vdd), .B(_1507__bF_buf7), );
  OAI21X1 OAI21X1_185 (.gnd(gnd), .A(_1505_), .Y(_320_), .vdd(vdd), .B(_1507__bF_buf6), .C(_1508_), );
  INVX2 INVX2_66 (.gnd(gnd), .A(regs_19__1_), .Y(_1509_), .vdd(vdd), );
  NAND2X1 NAND2X1_67 (.gnd(gnd), .A(wdata[1]), .Y(_1510_), .vdd(vdd), .B(_1507__bF_buf5), );
  OAI21X1 OAI21X1_186 (.gnd(gnd), .A(_1509_), .Y(_331_), .vdd(vdd), .B(_1507__bF_buf4), .C(_1510_), );
  INVX2 INVX2_67 (.gnd(gnd), .A(regs_19__2_), .Y(_1511_), .vdd(vdd), );
  NAND2X1 NAND2X1_68 (.gnd(gnd), .A(wdata[2]), .Y(_1512_), .vdd(vdd), .B(_1507__bF_buf3), );
  OAI21X1 OAI21X1_187 (.gnd(gnd), .A(_1511_), .Y(_342_), .vdd(vdd), .B(_1507__bF_buf2), .C(_1512_), );
  INVX2 INVX2_68 (.gnd(gnd), .A(regs_19__3_), .Y(_1513_), .vdd(vdd), );
  NAND2X1 NAND2X1_69 (.gnd(gnd), .A(wdata[3]), .Y(_1514_), .vdd(vdd), .B(_1507__bF_buf1), );
  OAI21X1 OAI21X1_188 (.gnd(gnd), .A(_1513_), .Y(_345_), .vdd(vdd), .B(_1507__bF_buf0), .C(_1514_), );
  INVX2 INVX2_69 (.gnd(gnd), .A(regs_19__4_), .Y(_1515_), .vdd(vdd), );
  NAND2X1 NAND2X1_70 (.gnd(gnd), .A(wdata[4]), .Y(_1516_), .vdd(vdd), .B(_1507__bF_buf7), );
  OAI21X1 OAI21X1_189 (.gnd(gnd), .A(_1515_), .Y(_346_), .vdd(vdd), .B(_1507__bF_buf6), .C(_1516_), );
  INVX2 INVX2_70 (.gnd(gnd), .A(regs_19__5_), .Y(_1517_), .vdd(vdd), );
  NAND2X1 NAND2X1_71 (.gnd(gnd), .A(wdata[5]), .Y(_1518_), .vdd(vdd), .B(_1507__bF_buf5), );
  OAI21X1 OAI21X1_190 (.gnd(gnd), .A(_1517_), .Y(_347_), .vdd(vdd), .B(_1507__bF_buf4), .C(_1518_), );
  INVX2 INVX2_71 (.gnd(gnd), .A(regs_19__6_), .Y(_1519_), .vdd(vdd), );
  NAND2X1 NAND2X1_72 (.gnd(gnd), .A(wdata[6]), .Y(_1520_), .vdd(vdd), .B(_1507__bF_buf3), );
  OAI21X1 OAI21X1_191 (.gnd(gnd), .A(_1519_), .Y(_348_), .vdd(vdd), .B(_1507__bF_buf2), .C(_1520_), );
  INVX2 INVX2_72 (.gnd(gnd), .A(regs_19__7_), .Y(_1521_), .vdd(vdd), );
  NAND2X1 NAND2X1_73 (.gnd(gnd), .A(wdata[7]), .Y(_1522_), .vdd(vdd), .B(_1507__bF_buf1), );
  OAI21X1 OAI21X1_192 (.gnd(gnd), .A(_1521_), .Y(_349_), .vdd(vdd), .B(_1507__bF_buf0), .C(_1522_), );
  INVX2 INVX2_73 (.gnd(gnd), .A(regs_19__8_), .Y(_1523_), .vdd(vdd), );
  NAND2X1 NAND2X1_74 (.gnd(gnd), .A(wdata[8]), .Y(_1524_), .vdd(vdd), .B(_1507__bF_buf7), );
  OAI21X1 OAI21X1_193 (.gnd(gnd), .A(_1523_), .Y(_350_), .vdd(vdd), .B(_1507__bF_buf6), .C(_1524_), );
  INVX2 INVX2_74 (.gnd(gnd), .A(regs_19__9_), .Y(_1525_), .vdd(vdd), );
  NAND2X1 NAND2X1_75 (.gnd(gnd), .A(wdata[9]), .Y(_1526_), .vdd(vdd), .B(_1507__bF_buf5), );
  OAI21X1 OAI21X1_194 (.gnd(gnd), .A(_1525_), .Y(_351_), .vdd(vdd), .B(_1507__bF_buf4), .C(_1526_), );
  INVX2 INVX2_75 (.gnd(gnd), .A(regs_19__10_), .Y(_1527_), .vdd(vdd), );
  NAND2X1 NAND2X1_76 (.gnd(gnd), .A(wdata[10]), .Y(_1528_), .vdd(vdd), .B(_1507__bF_buf3), );
  OAI21X1 OAI21X1_195 (.gnd(gnd), .A(_1527_), .Y(_321_), .vdd(vdd), .B(_1507__bF_buf2), .C(_1528_), );
  INVX2 INVX2_76 (.gnd(gnd), .A(regs_19__11_), .Y(_1529_), .vdd(vdd), );
  NAND2X1 NAND2X1_77 (.gnd(gnd), .A(wdata[11]), .Y(_1530_), .vdd(vdd), .B(_1507__bF_buf1), );
  OAI21X1 OAI21X1_196 (.gnd(gnd), .A(_1529_), .Y(_322_), .vdd(vdd), .B(_1507__bF_buf0), .C(_1530_), );
  INVX2 INVX2_77 (.gnd(gnd), .A(regs_19__12_), .Y(_1531_), .vdd(vdd), );
  NAND2X1 NAND2X1_78 (.gnd(gnd), .A(wdata[12]), .Y(_1532_), .vdd(vdd), .B(_1507__bF_buf7), );
  OAI21X1 OAI21X1_197 (.gnd(gnd), .A(_1531_), .Y(_323_), .vdd(vdd), .B(_1507__bF_buf6), .C(_1532_), );
  INVX2 INVX2_78 (.gnd(gnd), .A(regs_19__13_), .Y(_1533_), .vdd(vdd), );
  NAND2X1 NAND2X1_79 (.gnd(gnd), .A(wdata[13]), .Y(_1534_), .vdd(vdd), .B(_1507__bF_buf5), );
  OAI21X1 OAI21X1_198 (.gnd(gnd), .A(_1533_), .Y(_324_), .vdd(vdd), .B(_1507__bF_buf4), .C(_1534_), );
  INVX2 INVX2_79 (.gnd(gnd), .A(regs_19__14_), .Y(_1535_), .vdd(vdd), );
  NAND2X1 NAND2X1_80 (.gnd(gnd), .A(wdata[14]), .Y(_1536_), .vdd(vdd), .B(_1507__bF_buf3), );
  OAI21X1 OAI21X1_199 (.gnd(gnd), .A(_1535_), .Y(_325_), .vdd(vdd), .B(_1507__bF_buf2), .C(_1536_), );
  INVX2 INVX2_80 (.gnd(gnd), .A(regs_19__15_), .Y(_1537_), .vdd(vdd), );
  NAND2X1 NAND2X1_81 (.gnd(gnd), .A(wdata[15]), .Y(_1538_), .vdd(vdd), .B(_1507__bF_buf1), );
  OAI21X1 OAI21X1_200 (.gnd(gnd), .A(_1537_), .Y(_326_), .vdd(vdd), .B(_1507__bF_buf0), .C(_1538_), );
  INVX2 INVX2_81 (.gnd(gnd), .A(regs_19__16_), .Y(_1539_), .vdd(vdd), );
  NAND2X1 NAND2X1_82 (.gnd(gnd), .A(wdata[16]), .Y(_1540_), .vdd(vdd), .B(_1507__bF_buf7), );
  OAI21X1 OAI21X1_201 (.gnd(gnd), .A(_1539_), .Y(_327_), .vdd(vdd), .B(_1507__bF_buf6), .C(_1540_), );
  INVX2 INVX2_82 (.gnd(gnd), .A(regs_19__17_), .Y(_1541_), .vdd(vdd), );
  NAND2X1 NAND2X1_83 (.gnd(gnd), .A(wdata[17]), .Y(_1542_), .vdd(vdd), .B(_1507__bF_buf5), );
  OAI21X1 OAI21X1_202 (.gnd(gnd), .A(_1541_), .Y(_328_), .vdd(vdd), .B(_1507__bF_buf4), .C(_1542_), );
  INVX2 INVX2_83 (.gnd(gnd), .A(regs_19__18_), .Y(_1543_), .vdd(vdd), );
  NAND2X1 NAND2X1_84 (.gnd(gnd), .A(wdata[18]), .Y(_1544_), .vdd(vdd), .B(_1507__bF_buf3), );
  OAI21X1 OAI21X1_203 (.gnd(gnd), .A(_1543_), .Y(_329_), .vdd(vdd), .B(_1507__bF_buf2), .C(_1544_), );
  INVX2 INVX2_84 (.gnd(gnd), .A(regs_19__19_), .Y(_1545_), .vdd(vdd), );
  NAND2X1 NAND2X1_85 (.gnd(gnd), .A(wdata[19]), .Y(_1546_), .vdd(vdd), .B(_1507__bF_buf1), );
  OAI21X1 OAI21X1_204 (.gnd(gnd), .A(_1545_), .Y(_330_), .vdd(vdd), .B(_1507__bF_buf0), .C(_1546_), );
  INVX2 INVX2_85 (.gnd(gnd), .A(regs_19__20_), .Y(_1547_), .vdd(vdd), );
  NAND2X1 NAND2X1_86 (.gnd(gnd), .A(wdata[20]), .Y(_1548_), .vdd(vdd), .B(_1507__bF_buf7), );
  OAI21X1 OAI21X1_205 (.gnd(gnd), .A(_1547_), .Y(_332_), .vdd(vdd), .B(_1507__bF_buf6), .C(_1548_), );
  INVX2 INVX2_86 (.gnd(gnd), .A(regs_19__21_), .Y(_1549_), .vdd(vdd), );
  NAND2X1 NAND2X1_87 (.gnd(gnd), .A(wdata[21]), .Y(_1550_), .vdd(vdd), .B(_1507__bF_buf5), );
  OAI21X1 OAI21X1_206 (.gnd(gnd), .A(_1549_), .Y(_333_), .vdd(vdd), .B(_1507__bF_buf4), .C(_1550_), );
  INVX2 INVX2_87 (.gnd(gnd), .A(regs_19__22_), .Y(_1551_), .vdd(vdd), );
  NAND2X1 NAND2X1_88 (.gnd(gnd), .A(wdata[22]), .Y(_1552_), .vdd(vdd), .B(_1507__bF_buf3), );
  OAI21X1 OAI21X1_207 (.gnd(gnd), .A(_1551_), .Y(_334_), .vdd(vdd), .B(_1507__bF_buf2), .C(_1552_), );
  INVX2 INVX2_88 (.gnd(gnd), .A(regs_19__23_), .Y(_1553_), .vdd(vdd), );
  NAND2X1 NAND2X1_89 (.gnd(gnd), .A(wdata[23]), .Y(_1554_), .vdd(vdd), .B(_1507__bF_buf1), );
  OAI21X1 OAI21X1_208 (.gnd(gnd), .A(_1553_), .Y(_335_), .vdd(vdd), .B(_1507__bF_buf0), .C(_1554_), );
  INVX2 INVX2_89 (.gnd(gnd), .A(regs_19__24_), .Y(_1555_), .vdd(vdd), );
  NAND2X1 NAND2X1_90 (.gnd(gnd), .A(wdata[24]), .Y(_1556_), .vdd(vdd), .B(_1507__bF_buf7), );
  OAI21X1 OAI21X1_209 (.gnd(gnd), .A(_1555_), .Y(_336_), .vdd(vdd), .B(_1507__bF_buf6), .C(_1556_), );
  INVX2 INVX2_90 (.gnd(gnd), .A(regs_19__25_), .Y(_1557_), .vdd(vdd), );
  NAND2X1 NAND2X1_91 (.gnd(gnd), .A(wdata[25]), .Y(_1558_), .vdd(vdd), .B(_1507__bF_buf5), );
  OAI21X1 OAI21X1_210 (.gnd(gnd), .A(_1557_), .Y(_337_), .vdd(vdd), .B(_1507__bF_buf4), .C(_1558_), );
  INVX2 INVX2_91 (.gnd(gnd), .A(regs_19__26_), .Y(_1559_), .vdd(vdd), );
  NAND2X1 NAND2X1_92 (.gnd(gnd), .A(wdata[26]), .Y(_1560_), .vdd(vdd), .B(_1507__bF_buf3), );
  OAI21X1 OAI21X1_211 (.gnd(gnd), .A(_1559_), .Y(_338_), .vdd(vdd), .B(_1507__bF_buf2), .C(_1560_), );
  INVX2 INVX2_92 (.gnd(gnd), .A(regs_19__27_), .Y(_1561_), .vdd(vdd), );
  NAND2X1 NAND2X1_93 (.gnd(gnd), .A(wdata[27]), .Y(_1562_), .vdd(vdd), .B(_1507__bF_buf1), );
  OAI21X1 OAI21X1_212 (.gnd(gnd), .A(_1561_), .Y(_339_), .vdd(vdd), .B(_1507__bF_buf0), .C(_1562_), );
  INVX2 INVX2_93 (.gnd(gnd), .A(regs_19__28_), .Y(_1563_), .vdd(vdd), );
  NAND2X1 NAND2X1_94 (.gnd(gnd), .A(wdata[28]), .Y(_1564_), .vdd(vdd), .B(_1507__bF_buf7), );
  OAI21X1 OAI21X1_213 (.gnd(gnd), .A(_1563_), .Y(_340_), .vdd(vdd), .B(_1507__bF_buf6), .C(_1564_), );
  INVX2 INVX2_94 (.gnd(gnd), .A(regs_19__29_), .Y(_1565_), .vdd(vdd), );
  NAND2X1 NAND2X1_95 (.gnd(gnd), .A(wdata[29]), .Y(_1566_), .vdd(vdd), .B(_1507__bF_buf5), );
  OAI21X1 OAI21X1_214 (.gnd(gnd), .A(_1565_), .Y(_341_), .vdd(vdd), .B(_1507__bF_buf4), .C(_1566_), );
  INVX2 INVX2_95 (.gnd(gnd), .A(regs_19__30_), .Y(_1567_), .vdd(vdd), );
  NAND2X1 NAND2X1_96 (.gnd(gnd), .A(wdata[30]), .Y(_1568_), .vdd(vdd), .B(_1507__bF_buf3), );
  OAI21X1 OAI21X1_215 (.gnd(gnd), .A(_1567_), .Y(_343_), .vdd(vdd), .B(_1507__bF_buf2), .C(_1568_), );
  INVX2 INVX2_96 (.gnd(gnd), .A(regs_19__31_), .Y(_1569_), .vdd(vdd), );
  NAND2X1 NAND2X1_97 (.gnd(gnd), .A(wdata[31]), .Y(_1570_), .vdd(vdd), .B(_1507__bF_buf1), );
  OAI21X1 OAI21X1_216 (.gnd(gnd), .A(_1569_), .Y(_344_), .vdd(vdd), .B(_1507__bF_buf0), .C(_1570_), );
  NOR2X1 NOR2X1_37 (.gnd(gnd), .A(_1001__bF_buf8), .Y(_1571_), .vdd(vdd), .B(_1506__bF_buf4), );
  NOR2X1 NOR2X1_38 (.gnd(gnd), .A(regs_18__0_), .Y(_1572_), .vdd(vdd), .B(_1571__bF_buf7), );
  AOI21X1 AOI21X1_33 (.gnd(gnd), .A(_992__bF_buf1), .Y(_288_), .vdd(vdd), .B(_1571__bF_buf6), .C(_1572_), );
  NOR2X1 NOR2X1_39 (.gnd(gnd), .A(regs_18__1_), .Y(_1573_), .vdd(vdd), .B(_1571__bF_buf5), );
  AOI21X1 AOI21X1_34 (.gnd(gnd), .A(_1003__bF_buf1), .Y(_299_), .vdd(vdd), .B(_1571__bF_buf4), .C(_1573_), );
  NOR2X1 NOR2X1_40 (.gnd(gnd), .A(regs_18__2_), .Y(_1574_), .vdd(vdd), .B(_1571__bF_buf3), );
  AOI21X1 AOI21X1_35 (.gnd(gnd), .A(_1005__bF_buf1), .Y(_310_), .vdd(vdd), .B(_1571__bF_buf2), .C(_1574_), );
  NOR2X1 NOR2X1_41 (.gnd(gnd), .A(regs_18__3_), .Y(_1575_), .vdd(vdd), .B(_1571__bF_buf1), );
  AOI21X1 AOI21X1_36 (.gnd(gnd), .A(_1007__bF_buf1), .Y(_313_), .vdd(vdd), .B(_1571__bF_buf0), .C(_1575_), );
  NOR2X1 NOR2X1_42 (.gnd(gnd), .A(regs_18__4_), .Y(_1576_), .vdd(vdd), .B(_1571__bF_buf7), );
  AOI21X1 AOI21X1_37 (.gnd(gnd), .A(_1009__bF_buf0), .Y(_314_), .vdd(vdd), .B(_1571__bF_buf6), .C(_1576_), );
  NOR2X1 NOR2X1_43 (.gnd(gnd), .A(regs_18__5_), .Y(_1577_), .vdd(vdd), .B(_1571__bF_buf5), );
  AOI21X1 AOI21X1_38 (.gnd(gnd), .A(_1011__bF_buf0), .Y(_315_), .vdd(vdd), .B(_1571__bF_buf4), .C(_1577_), );
  NOR2X1 NOR2X1_44 (.gnd(gnd), .A(regs_18__6_), .Y(_1578_), .vdd(vdd), .B(_1571__bF_buf3), );
  AOI21X1 AOI21X1_39 (.gnd(gnd), .A(_1013__bF_buf0), .Y(_316_), .vdd(vdd), .B(_1571__bF_buf2), .C(_1578_), );
  NOR2X1 NOR2X1_45 (.gnd(gnd), .A(regs_18__7_), .Y(_1579_), .vdd(vdd), .B(_1571__bF_buf1), );
  AOI21X1 AOI21X1_40 (.gnd(gnd), .A(_1015__bF_buf0), .Y(_317_), .vdd(vdd), .B(_1571__bF_buf0), .C(_1579_), );
  NOR2X1 NOR2X1_46 (.gnd(gnd), .A(regs_18__8_), .Y(_1580_), .vdd(vdd), .B(_1571__bF_buf7), );
  AOI21X1 AOI21X1_41 (.gnd(gnd), .A(_1017__bF_buf0), .Y(_318_), .vdd(vdd), .B(_1571__bF_buf6), .C(_1580_), );
  NOR2X1 NOR2X1_47 (.gnd(gnd), .A(regs_18__9_), .Y(_1581_), .vdd(vdd), .B(_1571__bF_buf5), );
  AOI21X1 AOI21X1_42 (.gnd(gnd), .A(_1019__bF_buf0), .Y(_319_), .vdd(vdd), .B(_1571__bF_buf4), .C(_1581_), );
  NOR2X1 NOR2X1_48 (.gnd(gnd), .A(regs_18__10_), .Y(_1582_), .vdd(vdd), .B(_1571__bF_buf3), );
  AOI21X1 AOI21X1_43 (.gnd(gnd), .A(_1021__bF_buf0), .Y(_289_), .vdd(vdd), .B(_1571__bF_buf2), .C(_1582_), );
  NOR2X1 NOR2X1_49 (.gnd(gnd), .A(regs_18__11_), .Y(_1583_), .vdd(vdd), .B(_1571__bF_buf1), );
  AOI21X1 AOI21X1_44 (.gnd(gnd), .A(_1023__bF_buf0), .Y(_290_), .vdd(vdd), .B(_1571__bF_buf0), .C(_1583_), );
  NOR2X1 NOR2X1_50 (.gnd(gnd), .A(regs_18__12_), .Y(_1584_), .vdd(vdd), .B(_1571__bF_buf7), );
  AOI21X1 AOI21X1_45 (.gnd(gnd), .A(_1025__bF_buf0), .Y(_291_), .vdd(vdd), .B(_1571__bF_buf6), .C(_1584_), );
  NOR2X1 NOR2X1_51 (.gnd(gnd), .A(regs_18__13_), .Y(_1585_), .vdd(vdd), .B(_1571__bF_buf5), );
  AOI21X1 AOI21X1_46 (.gnd(gnd), .A(_1027__bF_buf0), .Y(_292_), .vdd(vdd), .B(_1571__bF_buf4), .C(_1585_), );
  NOR2X1 NOR2X1_52 (.gnd(gnd), .A(regs_18__14_), .Y(_1586_), .vdd(vdd), .B(_1571__bF_buf3), );
  AOI21X1 AOI21X1_47 (.gnd(gnd), .A(_1029__bF_buf0), .Y(_293_), .vdd(vdd), .B(_1571__bF_buf2), .C(_1586_), );
  NOR2X1 NOR2X1_53 (.gnd(gnd), .A(regs_18__15_), .Y(_1587_), .vdd(vdd), .B(_1571__bF_buf1), );
  AOI21X1 AOI21X1_48 (.gnd(gnd), .A(_1031__bF_buf0), .Y(_294_), .vdd(vdd), .B(_1571__bF_buf0), .C(_1587_), );
  NOR2X1 NOR2X1_54 (.gnd(gnd), .A(regs_18__16_), .Y(_1588_), .vdd(vdd), .B(_1571__bF_buf7), );
  AOI21X1 AOI21X1_49 (.gnd(gnd), .A(_1033__bF_buf0), .Y(_295_), .vdd(vdd), .B(_1571__bF_buf6), .C(_1588_), );
  NOR2X1 NOR2X1_55 (.gnd(gnd), .A(regs_18__17_), .Y(_1589_), .vdd(vdd), .B(_1571__bF_buf5), );
  AOI21X1 AOI21X1_50 (.gnd(gnd), .A(_1035__bF_buf0), .Y(_296_), .vdd(vdd), .B(_1571__bF_buf4), .C(_1589_), );
  NOR2X1 NOR2X1_56 (.gnd(gnd), .A(regs_18__18_), .Y(_1590_), .vdd(vdd), .B(_1571__bF_buf3), );
  AOI21X1 AOI21X1_51 (.gnd(gnd), .A(_1037__bF_buf0), .Y(_297_), .vdd(vdd), .B(_1571__bF_buf2), .C(_1590_), );
  NOR2X1 NOR2X1_57 (.gnd(gnd), .A(regs_18__19_), .Y(_1591_), .vdd(vdd), .B(_1571__bF_buf1), );
  AOI21X1 AOI21X1_52 (.gnd(gnd), .A(_1039__bF_buf0), .Y(_298_), .vdd(vdd), .B(_1571__bF_buf0), .C(_1591_), );
  NOR2X1 NOR2X1_58 (.gnd(gnd), .A(regs_18__20_), .Y(_1592_), .vdd(vdd), .B(_1571__bF_buf7), );
  AOI21X1 AOI21X1_53 (.gnd(gnd), .A(_1041__bF_buf0), .Y(_300_), .vdd(vdd), .B(_1571__bF_buf6), .C(_1592_), );
  NOR2X1 NOR2X1_59 (.gnd(gnd), .A(regs_18__21_), .Y(_1593_), .vdd(vdd), .B(_1571__bF_buf5), );
  AOI21X1 AOI21X1_54 (.gnd(gnd), .A(_1043__bF_buf0), .Y(_301_), .vdd(vdd), .B(_1571__bF_buf4), .C(_1593_), );
  NOR2X1 NOR2X1_60 (.gnd(gnd), .A(regs_18__22_), .Y(_1594_), .vdd(vdd), .B(_1571__bF_buf3), );
  AOI21X1 AOI21X1_55 (.gnd(gnd), .A(_1045__bF_buf0), .Y(_302_), .vdd(vdd), .B(_1571__bF_buf2), .C(_1594_), );
  NOR2X1 NOR2X1_61 (.gnd(gnd), .A(regs_18__23_), .Y(_1595_), .vdd(vdd), .B(_1571__bF_buf1), );
  AOI21X1 AOI21X1_56 (.gnd(gnd), .A(_1047__bF_buf0), .Y(_303_), .vdd(vdd), .B(_1571__bF_buf0), .C(_1595_), );
  NOR2X1 NOR2X1_62 (.gnd(gnd), .A(regs_18__24_), .Y(_1596_), .vdd(vdd), .B(_1571__bF_buf7), );
  AOI21X1 AOI21X1_57 (.gnd(gnd), .A(_1049__bF_buf0), .Y(_304_), .vdd(vdd), .B(_1571__bF_buf6), .C(_1596_), );
  NOR2X1 NOR2X1_63 (.gnd(gnd), .A(regs_18__25_), .Y(_1597_), .vdd(vdd), .B(_1571__bF_buf5), );
  AOI21X1 AOI21X1_58 (.gnd(gnd), .A(_1051__bF_buf0), .Y(_305_), .vdd(vdd), .B(_1571__bF_buf4), .C(_1597_), );
  NOR2X1 NOR2X1_64 (.gnd(gnd), .A(regs_18__26_), .Y(_1598_), .vdd(vdd), .B(_1571__bF_buf3), );
  AOI21X1 AOI21X1_59 (.gnd(gnd), .A(_1053__bF_buf0), .Y(_306_), .vdd(vdd), .B(_1571__bF_buf2), .C(_1598_), );
  NOR2X1 NOR2X1_65 (.gnd(gnd), .A(regs_18__27_), .Y(_1599_), .vdd(vdd), .B(_1571__bF_buf1), );
  AOI21X1 AOI21X1_60 (.gnd(gnd), .A(_1055__bF_buf0), .Y(_307_), .vdd(vdd), .B(_1571__bF_buf0), .C(_1599_), );
  NOR2X1 NOR2X1_66 (.gnd(gnd), .A(regs_18__28_), .Y(_1600_), .vdd(vdd), .B(_1571__bF_buf7), );
  AOI21X1 AOI21X1_61 (.gnd(gnd), .A(_1057__bF_buf0), .Y(_308_), .vdd(vdd), .B(_1571__bF_buf6), .C(_1600_), );
  NOR2X1 NOR2X1_67 (.gnd(gnd), .A(regs_18__29_), .Y(_1601_), .vdd(vdd), .B(_1571__bF_buf5), );
  AOI21X1 AOI21X1_62 (.gnd(gnd), .A(_1059__bF_buf0), .Y(_309_), .vdd(vdd), .B(_1571__bF_buf4), .C(_1601_), );
  NOR2X1 NOR2X1_68 (.gnd(gnd), .A(regs_18__30_), .Y(_1602_), .vdd(vdd), .B(_1571__bF_buf3), );
  AOI21X1 AOI21X1_63 (.gnd(gnd), .A(_1061__bF_buf0), .Y(_311_), .vdd(vdd), .B(_1571__bF_buf2), .C(_1602_), );
  NOR2X1 NOR2X1_69 (.gnd(gnd), .A(regs_18__31_), .Y(_1603_), .vdd(vdd), .B(_1571__bF_buf1), );
  AOI21X1 AOI21X1_64 (.gnd(gnd), .A(_1063__bF_buf0), .Y(_312_), .vdd(vdd), .B(_1571__bF_buf0), .C(_1603_), );
  INVX2 INVX2_97 (.gnd(gnd), .A(regs_17__0_), .Y(_1604_), .vdd(vdd), );
  NOR2X1 NOR2X1_70 (.gnd(gnd), .A(_1506__bF_buf3), .Y(_1605_), .vdd(vdd), .B(_1070__bF_buf9), );
  NAND2X1 NAND2X1_98 (.gnd(gnd), .A(wdata[0]), .Y(_1606_), .vdd(vdd), .B(_1605__bF_buf7), );
  OAI21X1 OAI21X1_217 (.gnd(gnd), .A(_1604_), .Y(_256_), .vdd(vdd), .B(_1605__bF_buf6), .C(_1606_), );
  INVX2 INVX2_98 (.gnd(gnd), .A(regs_17__1_), .Y(_1607_), .vdd(vdd), );
  NAND2X1 NAND2X1_99 (.gnd(gnd), .A(wdata[1]), .Y(_1608_), .vdd(vdd), .B(_1605__bF_buf5), );
  OAI21X1 OAI21X1_218 (.gnd(gnd), .A(_1607_), .Y(_267_), .vdd(vdd), .B(_1605__bF_buf4), .C(_1608_), );
  INVX2 INVX2_99 (.gnd(gnd), .A(regs_17__2_), .Y(_1609_), .vdd(vdd), );
  NAND2X1 NAND2X1_100 (.gnd(gnd), .A(wdata[2]), .Y(_1610_), .vdd(vdd), .B(_1605__bF_buf3), );
  OAI21X1 OAI21X1_219 (.gnd(gnd), .A(_1609_), .Y(_278_), .vdd(vdd), .B(_1605__bF_buf2), .C(_1610_), );
  INVX2 INVX2_100 (.gnd(gnd), .A(regs_17__3_), .Y(_1611_), .vdd(vdd), );
  NAND2X1 NAND2X1_101 (.gnd(gnd), .A(wdata[3]), .Y(_1612_), .vdd(vdd), .B(_1605__bF_buf1), );
  OAI21X1 OAI21X1_220 (.gnd(gnd), .A(_1611_), .Y(_281_), .vdd(vdd), .B(_1605__bF_buf0), .C(_1612_), );
  INVX2 INVX2_101 (.gnd(gnd), .A(regs_17__4_), .Y(_1613_), .vdd(vdd), );
  NAND2X1 NAND2X1_102 (.gnd(gnd), .A(wdata[4]), .Y(_1614_), .vdd(vdd), .B(_1605__bF_buf7), );
  OAI21X1 OAI21X1_221 (.gnd(gnd), .A(_1613_), .Y(_282_), .vdd(vdd), .B(_1605__bF_buf6), .C(_1614_), );
  INVX2 INVX2_102 (.gnd(gnd), .A(regs_17__5_), .Y(_1615_), .vdd(vdd), );
  NAND2X1 NAND2X1_103 (.gnd(gnd), .A(wdata[5]), .Y(_1616_), .vdd(vdd), .B(_1605__bF_buf5), );
  OAI21X1 OAI21X1_222 (.gnd(gnd), .A(_1615_), .Y(_283_), .vdd(vdd), .B(_1605__bF_buf4), .C(_1616_), );
  INVX2 INVX2_103 (.gnd(gnd), .A(regs_17__6_), .Y(_1617_), .vdd(vdd), );
  NAND2X1 NAND2X1_104 (.gnd(gnd), .A(wdata[6]), .Y(_1618_), .vdd(vdd), .B(_1605__bF_buf3), );
  OAI21X1 OAI21X1_223 (.gnd(gnd), .A(_1617_), .Y(_284_), .vdd(vdd), .B(_1605__bF_buf2), .C(_1618_), );
  INVX2 INVX2_104 (.gnd(gnd), .A(regs_17__7_), .Y(_1619_), .vdd(vdd), );
  NAND2X1 NAND2X1_105 (.gnd(gnd), .A(wdata[7]), .Y(_1620_), .vdd(vdd), .B(_1605__bF_buf1), );
  OAI21X1 OAI21X1_224 (.gnd(gnd), .A(_1619_), .Y(_285_), .vdd(vdd), .B(_1605__bF_buf0), .C(_1620_), );
  INVX2 INVX2_105 (.gnd(gnd), .A(regs_17__8_), .Y(_1621_), .vdd(vdd), );
  NAND2X1 NAND2X1_106 (.gnd(gnd), .A(wdata[8]), .Y(_1622_), .vdd(vdd), .B(_1605__bF_buf7), );
  OAI21X1 OAI21X1_225 (.gnd(gnd), .A(_1621_), .Y(_286_), .vdd(vdd), .B(_1605__bF_buf6), .C(_1622_), );
  INVX2 INVX2_106 (.gnd(gnd), .A(regs_17__9_), .Y(_1623_), .vdd(vdd), );
  NAND2X1 NAND2X1_107 (.gnd(gnd), .A(wdata[9]), .Y(_1624_), .vdd(vdd), .B(_1605__bF_buf5), );
  OAI21X1 OAI21X1_226 (.gnd(gnd), .A(_1623_), .Y(_287_), .vdd(vdd), .B(_1605__bF_buf4), .C(_1624_), );
  INVX2 INVX2_107 (.gnd(gnd), .A(regs_17__10_), .Y(_1625_), .vdd(vdd), );
  NAND2X1 NAND2X1_108 (.gnd(gnd), .A(wdata[10]), .Y(_1626_), .vdd(vdd), .B(_1605__bF_buf3), );
  OAI21X1 OAI21X1_227 (.gnd(gnd), .A(_1625_), .Y(_257_), .vdd(vdd), .B(_1605__bF_buf2), .C(_1626_), );
  INVX2 INVX2_108 (.gnd(gnd), .A(regs_17__11_), .Y(_1627_), .vdd(vdd), );
  NAND2X1 NAND2X1_109 (.gnd(gnd), .A(wdata[11]), .Y(_1628_), .vdd(vdd), .B(_1605__bF_buf1), );
  OAI21X1 OAI21X1_228 (.gnd(gnd), .A(_1627_), .Y(_258_), .vdd(vdd), .B(_1605__bF_buf0), .C(_1628_), );
  INVX2 INVX2_109 (.gnd(gnd), .A(regs_17__12_), .Y(_1629_), .vdd(vdd), );
  NAND2X1 NAND2X1_110 (.gnd(gnd), .A(wdata[12]), .Y(_1630_), .vdd(vdd), .B(_1605__bF_buf7), );
  OAI21X1 OAI21X1_229 (.gnd(gnd), .A(_1629_), .Y(_259_), .vdd(vdd), .B(_1605__bF_buf6), .C(_1630_), );
  INVX2 INVX2_110 (.gnd(gnd), .A(regs_17__13_), .Y(_1631_), .vdd(vdd), );
  NAND2X1 NAND2X1_111 (.gnd(gnd), .A(wdata[13]), .Y(_1632_), .vdd(vdd), .B(_1605__bF_buf5), );
  OAI21X1 OAI21X1_230 (.gnd(gnd), .A(_1631_), .Y(_260_), .vdd(vdd), .B(_1605__bF_buf4), .C(_1632_), );
  INVX2 INVX2_111 (.gnd(gnd), .A(regs_17__14_), .Y(_1633_), .vdd(vdd), );
  NAND2X1 NAND2X1_112 (.gnd(gnd), .A(wdata[14]), .Y(_1634_), .vdd(vdd), .B(_1605__bF_buf3), );
  OAI21X1 OAI21X1_231 (.gnd(gnd), .A(_1633_), .Y(_261_), .vdd(vdd), .B(_1605__bF_buf2), .C(_1634_), );
  INVX2 INVX2_112 (.gnd(gnd), .A(regs_17__15_), .Y(_1635_), .vdd(vdd), );
  NAND2X1 NAND2X1_113 (.gnd(gnd), .A(wdata[15]), .Y(_1636_), .vdd(vdd), .B(_1605__bF_buf1), );
  OAI21X1 OAI21X1_232 (.gnd(gnd), .A(_1635_), .Y(_262_), .vdd(vdd), .B(_1605__bF_buf0), .C(_1636_), );
  INVX2 INVX2_113 (.gnd(gnd), .A(regs_17__16_), .Y(_1637_), .vdd(vdd), );
  NAND2X1 NAND2X1_114 (.gnd(gnd), .A(wdata[16]), .Y(_1638_), .vdd(vdd), .B(_1605__bF_buf7), );
  OAI21X1 OAI21X1_233 (.gnd(gnd), .A(_1637_), .Y(_263_), .vdd(vdd), .B(_1605__bF_buf6), .C(_1638_), );
  INVX2 INVX2_114 (.gnd(gnd), .A(regs_17__17_), .Y(_1639_), .vdd(vdd), );
  NAND2X1 NAND2X1_115 (.gnd(gnd), .A(wdata[17]), .Y(_1640_), .vdd(vdd), .B(_1605__bF_buf5), );
  OAI21X1 OAI21X1_234 (.gnd(gnd), .A(_1639_), .Y(_264_), .vdd(vdd), .B(_1605__bF_buf4), .C(_1640_), );
  INVX2 INVX2_115 (.gnd(gnd), .A(regs_17__18_), .Y(_1641_), .vdd(vdd), );
  NAND2X1 NAND2X1_116 (.gnd(gnd), .A(wdata[18]), .Y(_1642_), .vdd(vdd), .B(_1605__bF_buf3), );
  OAI21X1 OAI21X1_235 (.gnd(gnd), .A(_1641_), .Y(_265_), .vdd(vdd), .B(_1605__bF_buf2), .C(_1642_), );
  INVX2 INVX2_116 (.gnd(gnd), .A(regs_17__19_), .Y(_1643_), .vdd(vdd), );
  NAND2X1 NAND2X1_117 (.gnd(gnd), .A(wdata[19]), .Y(_1644_), .vdd(vdd), .B(_1605__bF_buf1), );
  OAI21X1 OAI21X1_236 (.gnd(gnd), .A(_1643_), .Y(_266_), .vdd(vdd), .B(_1605__bF_buf0), .C(_1644_), );
  INVX2 INVX2_117 (.gnd(gnd), .A(regs_17__20_), .Y(_1645_), .vdd(vdd), );
  NAND2X1 NAND2X1_118 (.gnd(gnd), .A(wdata[20]), .Y(_1646_), .vdd(vdd), .B(_1605__bF_buf7), );
  OAI21X1 OAI21X1_237 (.gnd(gnd), .A(_1645_), .Y(_268_), .vdd(vdd), .B(_1605__bF_buf6), .C(_1646_), );
  INVX2 INVX2_118 (.gnd(gnd), .A(regs_17__21_), .Y(_1647_), .vdd(vdd), );
  NAND2X1 NAND2X1_119 (.gnd(gnd), .A(wdata[21]), .Y(_1648_), .vdd(vdd), .B(_1605__bF_buf5), );
  OAI21X1 OAI21X1_238 (.gnd(gnd), .A(_1647_), .Y(_269_), .vdd(vdd), .B(_1605__bF_buf4), .C(_1648_), );
  INVX2 INVX2_119 (.gnd(gnd), .A(regs_17__22_), .Y(_1649_), .vdd(vdd), );
  NAND2X1 NAND2X1_120 (.gnd(gnd), .A(wdata[22]), .Y(_1650_), .vdd(vdd), .B(_1605__bF_buf3), );
  OAI21X1 OAI21X1_239 (.gnd(gnd), .A(_1649_), .Y(_270_), .vdd(vdd), .B(_1605__bF_buf2), .C(_1650_), );
  INVX2 INVX2_120 (.gnd(gnd), .A(regs_17__23_), .Y(_1651_), .vdd(vdd), );
  NAND2X1 NAND2X1_121 (.gnd(gnd), .A(wdata[23]), .Y(_1652_), .vdd(vdd), .B(_1605__bF_buf1), );
  OAI21X1 OAI21X1_240 (.gnd(gnd), .A(_1651_), .Y(_271_), .vdd(vdd), .B(_1605__bF_buf0), .C(_1652_), );
  INVX2 INVX2_121 (.gnd(gnd), .A(regs_17__24_), .Y(_1653_), .vdd(vdd), );
  NAND2X1 NAND2X1_122 (.gnd(gnd), .A(wdata[24]), .Y(_1654_), .vdd(vdd), .B(_1605__bF_buf7), );
  OAI21X1 OAI21X1_241 (.gnd(gnd), .A(_1653_), .Y(_272_), .vdd(vdd), .B(_1605__bF_buf6), .C(_1654_), );
  INVX2 INVX2_122 (.gnd(gnd), .A(regs_17__25_), .Y(_1655_), .vdd(vdd), );
  NAND2X1 NAND2X1_123 (.gnd(gnd), .A(wdata[25]), .Y(_1656_), .vdd(vdd), .B(_1605__bF_buf5), );
  OAI21X1 OAI21X1_242 (.gnd(gnd), .A(_1655_), .Y(_273_), .vdd(vdd), .B(_1605__bF_buf4), .C(_1656_), );
  INVX2 INVX2_123 (.gnd(gnd), .A(regs_17__26_), .Y(_1657_), .vdd(vdd), );
  NAND2X1 NAND2X1_124 (.gnd(gnd), .A(wdata[26]), .Y(_1658_), .vdd(vdd), .B(_1605__bF_buf3), );
  OAI21X1 OAI21X1_243 (.gnd(gnd), .A(_1657_), .Y(_274_), .vdd(vdd), .B(_1605__bF_buf2), .C(_1658_), );
  INVX2 INVX2_124 (.gnd(gnd), .A(regs_17__27_), .Y(_1659_), .vdd(vdd), );
  NAND2X1 NAND2X1_125 (.gnd(gnd), .A(wdata[27]), .Y(_1660_), .vdd(vdd), .B(_1605__bF_buf1), );
  OAI21X1 OAI21X1_244 (.gnd(gnd), .A(_1659_), .Y(_275_), .vdd(vdd), .B(_1605__bF_buf0), .C(_1660_), );
  INVX2 INVX2_125 (.gnd(gnd), .A(regs_17__28_), .Y(_1661_), .vdd(vdd), );
  NAND2X1 NAND2X1_126 (.gnd(gnd), .A(wdata[28]), .Y(_1662_), .vdd(vdd), .B(_1605__bF_buf7), );
  OAI21X1 OAI21X1_245 (.gnd(gnd), .A(_1661_), .Y(_276_), .vdd(vdd), .B(_1605__bF_buf6), .C(_1662_), );
  INVX2 INVX2_126 (.gnd(gnd), .A(regs_17__29_), .Y(_1663_), .vdd(vdd), );
  NAND2X1 NAND2X1_127 (.gnd(gnd), .A(wdata[29]), .Y(_1664_), .vdd(vdd), .B(_1605__bF_buf5), );
  OAI21X1 OAI21X1_246 (.gnd(gnd), .A(_1663_), .Y(_277_), .vdd(vdd), .B(_1605__bF_buf4), .C(_1664_), );
  INVX2 INVX2_127 (.gnd(gnd), .A(regs_17__30_), .Y(_1665_), .vdd(vdd), );
  NAND2X1 NAND2X1_128 (.gnd(gnd), .A(wdata[30]), .Y(_1666_), .vdd(vdd), .B(_1605__bF_buf3), );
  OAI21X1 OAI21X1_247 (.gnd(gnd), .A(_1665_), .Y(_279_), .vdd(vdd), .B(_1605__bF_buf2), .C(_1666_), );
  INVX2 INVX2_128 (.gnd(gnd), .A(regs_17__31_), .Y(_1667_), .vdd(vdd), );
  NAND2X1 NAND2X1_129 (.gnd(gnd), .A(wdata[31]), .Y(_1668_), .vdd(vdd), .B(_1605__bF_buf1), );
  OAI21X1 OAI21X1_248 (.gnd(gnd), .A(_1667_), .Y(_280_), .vdd(vdd), .B(_1605__bF_buf0), .C(_1668_), );
  OR2X2 OR2X2_4 (.gnd(gnd), .A(_1506__bF_buf2), .Y(_1669_), .vdd(vdd), .B(_1104__bF_buf13), );
  OAI21X1 OAI21X1_249 (.gnd(gnd), .A(_1506__bF_buf1), .Y(_1670_), .vdd(vdd), .B(_1104__bF_buf12), .C(regs_16__0_), );
  OAI21X1 OAI21X1_250 (.gnd(gnd), .A(_1669__bF_buf4), .Y(_224_), .vdd(vdd), .B(_992__bF_buf0), .C(_1670_), );
  OAI21X1 OAI21X1_251 (.gnd(gnd), .A(_1506__bF_buf0), .Y(_1671_), .vdd(vdd), .B(_1104__bF_buf11), .C(regs_16__1_), );
  OAI21X1 OAI21X1_252 (.gnd(gnd), .A(_1669__bF_buf3), .Y(_235_), .vdd(vdd), .B(_1003__bF_buf0), .C(_1671_), );
  OAI21X1 OAI21X1_253 (.gnd(gnd), .A(_1506__bF_buf5), .Y(_1672_), .vdd(vdd), .B(_1104__bF_buf10), .C(regs_16__2_), );
  OAI21X1 OAI21X1_254 (.gnd(gnd), .A(_1669__bF_buf2), .Y(_246_), .vdd(vdd), .B(_1005__bF_buf0), .C(_1672_), );
  OAI21X1 OAI21X1_255 (.gnd(gnd), .A(_1506__bF_buf4), .Y(_1673_), .vdd(vdd), .B(_1104__bF_buf9), .C(regs_16__3_), );
  OAI21X1 OAI21X1_256 (.gnd(gnd), .A(_1669__bF_buf1), .Y(_249_), .vdd(vdd), .B(_1007__bF_buf0), .C(_1673_), );
  OAI21X1 OAI21X1_257 (.gnd(gnd), .A(_1506__bF_buf3), .Y(_1674_), .vdd(vdd), .B(_1104__bF_buf8), .C(regs_16__4_), );
  OAI21X1 OAI21X1_258 (.gnd(gnd), .A(_1669__bF_buf0), .Y(_250_), .vdd(vdd), .B(_1009__bF_buf3), .C(_1674_), );
  OAI21X1 OAI21X1_259 (.gnd(gnd), .A(_1506__bF_buf2), .Y(_1675_), .vdd(vdd), .B(_1104__bF_buf7), .C(regs_16__5_), );
  OAI21X1 OAI21X1_260 (.gnd(gnd), .A(_1669__bF_buf4), .Y(_251_), .vdd(vdd), .B(_1011__bF_buf3), .C(_1675_), );
  OAI21X1 OAI21X1_261 (.gnd(gnd), .A(_1506__bF_buf1), .Y(_1676_), .vdd(vdd), .B(_1104__bF_buf6), .C(regs_16__6_), );
  OAI21X1 OAI21X1_262 (.gnd(gnd), .A(_1669__bF_buf3), .Y(_252_), .vdd(vdd), .B(_1013__bF_buf3), .C(_1676_), );
  OAI21X1 OAI21X1_263 (.gnd(gnd), .A(_1506__bF_buf0), .Y(_1677_), .vdd(vdd), .B(_1104__bF_buf5), .C(regs_16__7_), );
  OAI21X1 OAI21X1_264 (.gnd(gnd), .A(_1669__bF_buf2), .Y(_253_), .vdd(vdd), .B(_1015__bF_buf3), .C(_1677_), );
  OAI21X1 OAI21X1_265 (.gnd(gnd), .A(_1506__bF_buf5), .Y(_1678_), .vdd(vdd), .B(_1104__bF_buf4), .C(regs_16__8_), );
  OAI21X1 OAI21X1_266 (.gnd(gnd), .A(_1669__bF_buf1), .Y(_254_), .vdd(vdd), .B(_1017__bF_buf3), .C(_1678_), );
  OAI21X1 OAI21X1_267 (.gnd(gnd), .A(_1506__bF_buf4), .Y(_1679_), .vdd(vdd), .B(_1104__bF_buf3), .C(regs_16__9_), );
  OAI21X1 OAI21X1_268 (.gnd(gnd), .A(_1669__bF_buf0), .Y(_255_), .vdd(vdd), .B(_1019__bF_buf3), .C(_1679_), );
  OAI21X1 OAI21X1_269 (.gnd(gnd), .A(_1506__bF_buf3), .Y(_1680_), .vdd(vdd), .B(_1104__bF_buf2), .C(regs_16__10_), );
  OAI21X1 OAI21X1_270 (.gnd(gnd), .A(_1669__bF_buf4), .Y(_225_), .vdd(vdd), .B(_1021__bF_buf3), .C(_1680_), );
  OAI21X1 OAI21X1_271 (.gnd(gnd), .A(_1506__bF_buf2), .Y(_1681_), .vdd(vdd), .B(_1104__bF_buf1), .C(regs_16__11_), );
  OAI21X1 OAI21X1_272 (.gnd(gnd), .A(_1669__bF_buf3), .Y(_226_), .vdd(vdd), .B(_1023__bF_buf3), .C(_1681_), );
  OAI21X1 OAI21X1_273 (.gnd(gnd), .A(_1506__bF_buf1), .Y(_1682_), .vdd(vdd), .B(_1104__bF_buf0), .C(regs_16__12_), );
  OAI21X1 OAI21X1_274 (.gnd(gnd), .A(_1669__bF_buf2), .Y(_227_), .vdd(vdd), .B(_1025__bF_buf3), .C(_1682_), );
  OAI21X1 OAI21X1_275 (.gnd(gnd), .A(_1506__bF_buf0), .Y(_1683_), .vdd(vdd), .B(_1104__bF_buf14), .C(regs_16__13_), );
  OAI21X1 OAI21X1_276 (.gnd(gnd), .A(_1669__bF_buf1), .Y(_228_), .vdd(vdd), .B(_1027__bF_buf3), .C(_1683_), );
  OAI21X1 OAI21X1_277 (.gnd(gnd), .A(_1506__bF_buf5), .Y(_1684_), .vdd(vdd), .B(_1104__bF_buf13), .C(regs_16__14_), );
  OAI21X1 OAI21X1_278 (.gnd(gnd), .A(_1669__bF_buf0), .Y(_229_), .vdd(vdd), .B(_1029__bF_buf3), .C(_1684_), );
  OAI21X1 OAI21X1_279 (.gnd(gnd), .A(_1506__bF_buf4), .Y(_1685_), .vdd(vdd), .B(_1104__bF_buf12), .C(regs_16__15_), );
  OAI21X1 OAI21X1_280 (.gnd(gnd), .A(_1669__bF_buf4), .Y(_230_), .vdd(vdd), .B(_1031__bF_buf3), .C(_1685_), );
  OAI21X1 OAI21X1_281 (.gnd(gnd), .A(_1506__bF_buf3), .Y(_1686_), .vdd(vdd), .B(_1104__bF_buf11), .C(regs_16__16_), );
  OAI21X1 OAI21X1_282 (.gnd(gnd), .A(_1669__bF_buf3), .Y(_231_), .vdd(vdd), .B(_1033__bF_buf3), .C(_1686_), );
  OAI21X1 OAI21X1_283 (.gnd(gnd), .A(_1506__bF_buf2), .Y(_1687_), .vdd(vdd), .B(_1104__bF_buf10), .C(regs_16__17_), );
  OAI21X1 OAI21X1_284 (.gnd(gnd), .A(_1669__bF_buf2), .Y(_232_), .vdd(vdd), .B(_1035__bF_buf3), .C(_1687_), );
  OAI21X1 OAI21X1_285 (.gnd(gnd), .A(_1506__bF_buf1), .Y(_1688_), .vdd(vdd), .B(_1104__bF_buf9), .C(regs_16__18_), );
  OAI21X1 OAI21X1_286 (.gnd(gnd), .A(_1669__bF_buf1), .Y(_233_), .vdd(vdd), .B(_1037__bF_buf3), .C(_1688_), );
  OAI21X1 OAI21X1_287 (.gnd(gnd), .A(_1506__bF_buf0), .Y(_1689_), .vdd(vdd), .B(_1104__bF_buf8), .C(regs_16__19_), );
  OAI21X1 OAI21X1_288 (.gnd(gnd), .A(_1669__bF_buf0), .Y(_234_), .vdd(vdd), .B(_1039__bF_buf3), .C(_1689_), );
  OAI21X1 OAI21X1_289 (.gnd(gnd), .A(_1506__bF_buf5), .Y(_1690_), .vdd(vdd), .B(_1104__bF_buf7), .C(regs_16__20_), );
  OAI21X1 OAI21X1_290 (.gnd(gnd), .A(_1669__bF_buf4), .Y(_236_), .vdd(vdd), .B(_1041__bF_buf3), .C(_1690_), );
  OAI21X1 OAI21X1_291 (.gnd(gnd), .A(_1506__bF_buf4), .Y(_1691_), .vdd(vdd), .B(_1104__bF_buf6), .C(regs_16__21_), );
  OAI21X1 OAI21X1_292 (.gnd(gnd), .A(_1669__bF_buf3), .Y(_237_), .vdd(vdd), .B(_1043__bF_buf3), .C(_1691_), );
  OAI21X1 OAI21X1_293 (.gnd(gnd), .A(_1506__bF_buf3), .Y(_1692_), .vdd(vdd), .B(_1104__bF_buf5), .C(regs_16__22_), );
  OAI21X1 OAI21X1_294 (.gnd(gnd), .A(_1669__bF_buf2), .Y(_238_), .vdd(vdd), .B(_1045__bF_buf3), .C(_1692_), );
  OAI21X1 OAI21X1_295 (.gnd(gnd), .A(_1506__bF_buf2), .Y(_1693_), .vdd(vdd), .B(_1104__bF_buf4), .C(regs_16__23_), );
  OAI21X1 OAI21X1_296 (.gnd(gnd), .A(_1669__bF_buf1), .Y(_239_), .vdd(vdd), .B(_1047__bF_buf3), .C(_1693_), );
  OAI21X1 OAI21X1_297 (.gnd(gnd), .A(_1506__bF_buf1), .Y(_1694_), .vdd(vdd), .B(_1104__bF_buf3), .C(regs_16__24_), );
  OAI21X1 OAI21X1_298 (.gnd(gnd), .A(_1669__bF_buf0), .Y(_240_), .vdd(vdd), .B(_1049__bF_buf3), .C(_1694_), );
  OAI21X1 OAI21X1_299 (.gnd(gnd), .A(_1506__bF_buf0), .Y(_1695_), .vdd(vdd), .B(_1104__bF_buf2), .C(regs_16__25_), );
  OAI21X1 OAI21X1_300 (.gnd(gnd), .A(_1669__bF_buf4), .Y(_241_), .vdd(vdd), .B(_1051__bF_buf3), .C(_1695_), );
  OAI21X1 OAI21X1_301 (.gnd(gnd), .A(_1506__bF_buf5), .Y(_1696_), .vdd(vdd), .B(_1104__bF_buf1), .C(regs_16__26_), );
  OAI21X1 OAI21X1_302 (.Y(_242_), .A(_1669__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1053__bF_buf3), .C(_1696_), );
  OAI21X1 OAI21X1_303 (.Y(_1697_), .A(_1506__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf0), .C(regs_16__27_), );
  OAI21X1 OAI21X1_304 (.Y(_243_), .A(_1669__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1055__bF_buf3), .C(_1697_), );
  OAI21X1 OAI21X1_305 (.Y(_1698_), .A(_1506__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf14), .C(regs_16__28_), );
  OAI21X1 OAI21X1_306 (.Y(_244_), .A(_1669__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1057__bF_buf3), .C(_1698_), );
  OAI21X1 OAI21X1_307 (.Y(_1699_), .A(_1506__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf13), .C(regs_16__29_), );
  OAI21X1 OAI21X1_308 (.Y(_245_), .A(_1669__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1059__bF_buf3), .C(_1699_), );
  OAI21X1 OAI21X1_309 (.Y(_1700_), .A(_1506__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf12), .C(regs_16__30_), );
  OAI21X1 OAI21X1_310 (.Y(_247_), .A(_1669__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1061__bF_buf3), .C(_1700_), );
  OAI21X1 OAI21X1_311 (.Y(_1701_), .A(_1506__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf11), .C(regs_16__31_), );
  OAI21X1 OAI21X1_312 (.Y(_248_), .A(_1669__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1063__bF_buf3), .C(_1701_), );
  INVX2 INVX2_129 (.Y(_1702_), .A(regs_15__0_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_130 (.Y(_1703_), .A(waddr[4]), .gnd(gnd), .vdd(vdd), .B(_994_), );
  OR2X2 OR2X2_5 (.Y(_1704_), .A(_1703_), .gnd(gnd), .vdd(vdd), .B(waddr[2]), );
  NOR2X1 NOR2X1_71 (.Y(_1705_), .A(_1142__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1704__bF_buf5), );
  NAND2X1 NAND2X1_131 (.Y(_1706_), .A(wdata[0]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf7), );
  OAI21X1 OAI21X1_313 (.Y(_192_), .A(_1702_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf6), .C(_1706_), );
  INVX2 INVX2_130 (.Y(_1707_), .A(regs_15__1_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_132 (.Y(_1708_), .A(wdata[1]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf5), );
  OAI21X1 OAI21X1_314 (.Y(_203_), .A(_1707_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf4), .C(_1708_), );
  INVX2 INVX2_131 (.Y(_1709_), .A(regs_15__2_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_133 (.Y(_1710_), .A(wdata[2]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf3), );
  OAI21X1 OAI21X1_315 (.Y(_214_), .A(_1709_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf2), .C(_1710_), );
  INVX2 INVX2_132 (.Y(_1711_), .A(regs_15__3_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_134 (.Y(_1712_), .A(wdata[3]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf1), );
  OAI21X1 OAI21X1_316 (.Y(_217_), .A(_1711_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf0), .C(_1712_), );
  INVX2 INVX2_133 (.Y(_1713_), .A(regs_15__4_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_135 (.Y(_1714_), .A(wdata[4]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf7), );
  OAI21X1 OAI21X1_317 (.Y(_218_), .A(_1713_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf6), .C(_1714_), );
  INVX2 INVX2_134 (.Y(_1715_), .A(regs_15__5_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_136 (.Y(_1716_), .A(wdata[5]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf5), );
  OAI21X1 OAI21X1_318 (.Y(_219_), .A(_1715_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf4), .C(_1716_), );
  INVX2 INVX2_135 (.Y(_1717_), .A(regs_15__6_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_137 (.Y(_1718_), .A(wdata[6]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf3), );
  OAI21X1 OAI21X1_319 (.Y(_220_), .A(_1717_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf2), .C(_1718_), );
  INVX2 INVX2_136 (.Y(_1719_), .A(regs_15__7_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_138 (.Y(_1720_), .A(wdata[7]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf1), );
  OAI21X1 OAI21X1_320 (.Y(_221_), .A(_1719_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf0), .C(_1720_), );
  INVX2 INVX2_137 (.Y(_1721_), .A(regs_15__8_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_139 (.Y(_1722_), .A(wdata[8]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf7), );
  OAI21X1 OAI21X1_321 (.Y(_222_), .A(_1721_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf6), .C(_1722_), );
  INVX2 INVX2_138 (.Y(_1723_), .A(regs_15__9_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_140 (.Y(_1724_), .A(wdata[9]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf5), );
  OAI21X1 OAI21X1_322 (.Y(_223_), .A(_1723_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf4), .C(_1724_), );
  INVX2 INVX2_139 (.Y(_1725_), .A(regs_15__10_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_141 (.Y(_1726_), .A(wdata[10]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf3), );
  OAI21X1 OAI21X1_323 (.Y(_193_), .A(_1725_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf2), .C(_1726_), );
  INVX2 INVX2_140 (.Y(_1727_), .A(regs_15__11_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_142 (.Y(_1728_), .A(wdata[11]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf1), );
  OAI21X1 OAI21X1_324 (.Y(_194_), .A(_1727_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf0), .C(_1728_), );
  INVX2 INVX2_141 (.Y(_1729_), .A(regs_15__12_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_143 (.Y(_1730_), .A(wdata[12]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf7), );
  OAI21X1 OAI21X1_325 (.Y(_195_), .A(_1729_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf6), .C(_1730_), );
  INVX2 INVX2_142 (.Y(_1731_), .A(regs_15__13_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_144 (.Y(_1732_), .A(wdata[13]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf5), );
  OAI21X1 OAI21X1_326 (.Y(_196_), .A(_1731_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf4), .C(_1732_), );
  INVX2 INVX2_143 (.Y(_1733_), .A(regs_15__14_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_145 (.Y(_1734_), .A(wdata[14]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf3), );
  OAI21X1 OAI21X1_327 (.Y(_197_), .A(_1733_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf2), .C(_1734_), );
  INVX2 INVX2_144 (.Y(_1735_), .A(regs_15__15_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_146 (.Y(_1736_), .A(wdata[15]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf1), );
  OAI21X1 OAI21X1_328 (.Y(_198_), .A(_1735_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf0), .C(_1736_), );
  INVX2 INVX2_145 (.Y(_1737_), .A(regs_15__16_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_147 (.Y(_1738_), .A(wdata[16]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf7), );
  OAI21X1 OAI21X1_329 (.Y(_199_), .A(_1737_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf6), .C(_1738_), );
  INVX2 INVX2_146 (.Y(_1739_), .A(regs_15__17_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_148 (.Y(_1740_), .A(wdata[17]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf5), );
  OAI21X1 OAI21X1_330 (.Y(_200_), .A(_1739_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf4), .C(_1740_), );
  INVX2 INVX2_147 (.Y(_1741_), .A(regs_15__18_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_149 (.Y(_1742_), .A(wdata[18]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf3), );
  OAI21X1 OAI21X1_331 (.Y(_201_), .A(_1741_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf2), .C(_1742_), );
  INVX2 INVX2_148 (.Y(_1743_), .A(regs_15__19_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_150 (.Y(_1744_), .A(wdata[19]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf1), );
  OAI21X1 OAI21X1_332 (.Y(_202_), .A(_1743_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf0), .C(_1744_), );
  INVX2 INVX2_149 (.Y(_1745_), .A(regs_15__20_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_151 (.Y(_1746_), .A(wdata[20]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf7), );
  OAI21X1 OAI21X1_333 (.Y(_204_), .A(_1745_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf6), .C(_1746_), );
  INVX2 INVX2_150 (.Y(_1747_), .A(regs_15__21_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_152 (.Y(_1748_), .A(wdata[21]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf5), );
  OAI21X1 OAI21X1_334 (.Y(_205_), .A(_1747_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf4), .C(_1748_), );
  INVX2 INVX2_151 (.Y(_1749_), .A(regs_15__22_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_153 (.Y(_1750_), .A(wdata[22]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf3), );
  OAI21X1 OAI21X1_335 (.Y(_206_), .A(_1749_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf2), .C(_1750_), );
  INVX2 INVX2_152 (.Y(_1751_), .A(regs_15__23_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_154 (.Y(_1752_), .A(wdata[23]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf1), );
  OAI21X1 OAI21X1_336 (.Y(_207_), .A(_1751_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf0), .C(_1752_), );
  INVX2 INVX2_153 (.Y(_1753_), .A(regs_15__24_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_155 (.Y(_1754_), .A(wdata[24]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf7), );
  OAI21X1 OAI21X1_337 (.Y(_208_), .A(_1753_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf6), .C(_1754_), );
  INVX2 INVX2_154 (.Y(_1755_), .A(regs_15__25_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_156 (.Y(_1756_), .A(wdata[25]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf5), );
  OAI21X1 OAI21X1_338 (.Y(_209_), .A(_1755_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf4), .C(_1756_), );
  INVX2 INVX2_155 (.Y(_1757_), .A(regs_15__26_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_157 (.Y(_1758_), .A(wdata[26]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf3), );
  OAI21X1 OAI21X1_339 (.Y(_210_), .A(_1757_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf2), .C(_1758_), );
  INVX2 INVX2_156 (.Y(_1759_), .A(regs_15__27_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_158 (.Y(_1760_), .A(wdata[27]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf1), );
  OAI21X1 OAI21X1_340 (.Y(_211_), .A(_1759_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf0), .C(_1760_), );
  INVX2 INVX2_157 (.Y(_1761_), .A(regs_15__28_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_159 (.Y(_1762_), .A(wdata[28]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf7), );
  OAI21X1 OAI21X1_341 (.Y(_212_), .A(_1761_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf6), .C(_1762_), );
  INVX2 INVX2_158 (.Y(_1763_), .A(regs_15__29_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_160 (.Y(_1764_), .A(wdata[29]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf5), );
  OAI21X1 OAI21X1_342 (.Y(_213_), .A(_1763_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf4), .C(_1764_), );
  INVX2 INVX2_159 (.Y(_1765_), .A(regs_15__30_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_161 (.Y(_1766_), .A(wdata[30]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf3), );
  OAI21X1 OAI21X1_343 (.Y(_215_), .A(_1765_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf2), .C(_1766_), );
  INVX2 INVX2_160 (.Y(_1767_), .A(regs_15__31_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_162 (.Y(_1768_), .A(wdata[31]), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf1), );
  OAI21X1 OAI21X1_344 (.Y(_216_), .A(_1767_), .gnd(gnd), .vdd(vdd), .B(_1705__bF_buf0), .C(_1768_), );
  NOR2X1 NOR2X1_72 (.Y(_1769_), .A(_1001__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_1704__bF_buf4), );
  NOR2X1 NOR2X1_73 (.Y(_1770_), .A(regs_14__0_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf7), );
  AOI21X1 AOI21X1_65 (.Y(_160_), .A(_992__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf6), .C(_1770_), );
  NOR2X1 NOR2X1_74 (.Y(_1771_), .A(regs_14__1_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf5), );
  AOI21X1 AOI21X1_66 (.Y(_171_), .A(_1003__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf4), .C(_1771_), );
  NOR2X1 NOR2X1_75 (.Y(_1772_), .A(regs_14__2_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf3), );
  AOI21X1 AOI21X1_67 (.Y(_182_), .A(_1005__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf2), .C(_1772_), );
  NOR2X1 NOR2X1_76 (.Y(_1773_), .A(regs_14__3_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf1), );
  AOI21X1 AOI21X1_68 (.Y(_185_), .A(_1007__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf0), .C(_1773_), );
  NOR2X1 NOR2X1_77 (.Y(_1774_), .A(regs_14__4_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf7), );
  AOI21X1 AOI21X1_69 (.Y(_186_), .A(_1009__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf6), .C(_1774_), );
  NOR2X1 NOR2X1_78 (.Y(_1775_), .A(regs_14__5_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf5), );
  AOI21X1 AOI21X1_70 (.Y(_187_), .A(_1011__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf4), .C(_1775_), );
  NOR2X1 NOR2X1_79 (.Y(_1776_), .A(regs_14__6_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf3), );
  AOI21X1 AOI21X1_71 (.Y(_188_), .A(_1013__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf2), .C(_1776_), );
  NOR2X1 NOR2X1_80 (.Y(_1777_), .A(regs_14__7_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf1), );
  AOI21X1 AOI21X1_72 (.Y(_189_), .A(_1015__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf0), .C(_1777_), );
  NOR2X1 NOR2X1_81 (.Y(_1778_), .A(regs_14__8_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf7), );
  AOI21X1 AOI21X1_73 (.Y(_190_), .A(_1017__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf6), .C(_1778_), );
  NOR2X1 NOR2X1_82 (.Y(_1779_), .A(regs_14__9_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf5), );
  AOI21X1 AOI21X1_74 (.Y(_191_), .A(_1019__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf4), .C(_1779_), );
  NOR2X1 NOR2X1_83 (.Y(_1780_), .A(regs_14__10_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf3), );
  AOI21X1 AOI21X1_75 (.Y(_161_), .A(_1021__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf2), .C(_1780_), );
  NOR2X1 NOR2X1_84 (.Y(_1781_), .A(regs_14__11_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf1), );
  AOI21X1 AOI21X1_76 (.Y(_162_), .A(_1023__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf0), .C(_1781_), );
  NOR2X1 NOR2X1_85 (.Y(_1782_), .A(regs_14__12_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf7), );
  AOI21X1 AOI21X1_77 (.Y(_163_), .A(_1025__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf6), .C(_1782_), );
  NOR2X1 NOR2X1_86 (.Y(_1783_), .A(regs_14__13_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf5), );
  AOI21X1 AOI21X1_78 (.Y(_164_), .A(_1027__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf4), .C(_1783_), );
  NOR2X1 NOR2X1_87 (.Y(_1784_), .A(regs_14__14_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf3), );
  AOI21X1 AOI21X1_79 (.Y(_165_), .A(_1029__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf2), .C(_1784_), );
  NOR2X1 NOR2X1_88 (.Y(_1785_), .A(regs_14__15_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf1), );
  AOI21X1 AOI21X1_80 (.Y(_166_), .A(_1031__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf0), .C(_1785_), );
  NOR2X1 NOR2X1_89 (.Y(_1786_), .A(regs_14__16_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf7), );
  AOI21X1 AOI21X1_81 (.Y(_167_), .A(_1033__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf6), .C(_1786_), );
  NOR2X1 NOR2X1_90 (.Y(_1787_), .A(regs_14__17_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf5), );
  AOI21X1 AOI21X1_82 (.Y(_168_), .A(_1035__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf4), .C(_1787_), );
  NOR2X1 NOR2X1_91 (.Y(_1788_), .A(regs_14__18_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf3), );
  AOI21X1 AOI21X1_83 (.Y(_169_), .A(_1037__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf2), .C(_1788_), );
  NOR2X1 NOR2X1_92 (.Y(_1789_), .A(regs_14__19_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf1), );
  AOI21X1 AOI21X1_84 (.Y(_170_), .A(_1039__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf0), .C(_1789_), );
  NOR2X1 NOR2X1_93 (.Y(_1790_), .A(regs_14__20_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf7), );
  AOI21X1 AOI21X1_85 (.Y(_172_), .A(_1041__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf6), .C(_1790_), );
  NOR2X1 NOR2X1_94 (.Y(_1791_), .A(regs_14__21_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf5), );
  AOI21X1 AOI21X1_86 (.Y(_173_), .A(_1043__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf4), .C(_1791_), );
  NOR2X1 NOR2X1_95 (.Y(_1792_), .A(regs_14__22_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf3), );
  AOI21X1 AOI21X1_87 (.Y(_174_), .A(_1045__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf2), .C(_1792_), );
  NOR2X1 NOR2X1_96 (.Y(_1793_), .A(regs_14__23_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf1), );
  AOI21X1 AOI21X1_88 (.Y(_175_), .A(_1047__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf0), .C(_1793_), );
  NOR2X1 NOR2X1_97 (.Y(_1794_), .A(regs_14__24_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf7), );
  AOI21X1 AOI21X1_89 (.Y(_176_), .A(_1049__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf6), .C(_1794_), );
  NOR2X1 NOR2X1_98 (.Y(_1795_), .A(regs_14__25_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf5), );
  AOI21X1 AOI21X1_90 (.Y(_177_), .A(_1051__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf4), .C(_1795_), );
  NOR2X1 NOR2X1_99 (.Y(_1796_), .A(regs_14__26_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf3), );
  AOI21X1 AOI21X1_91 (.Y(_178_), .A(_1053__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf2), .C(_1796_), );
  NOR2X1 NOR2X1_100 (.Y(_1797_), .A(regs_14__27_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf1), );
  AOI21X1 AOI21X1_92 (.Y(_179_), .A(_1055__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf0), .C(_1797_), );
  NOR2X1 NOR2X1_101 (.Y(_1798_), .A(regs_14__28_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf7), );
  AOI21X1 AOI21X1_93 (.Y(_180_), .A(_1057__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf6), .C(_1798_), );
  NOR2X1 NOR2X1_102 (.Y(_1799_), .A(regs_14__29_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf5), );
  AOI21X1 AOI21X1_94 (.Y(_181_), .A(_1059__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf4), .C(_1799_), );
  NOR2X1 NOR2X1_103 (.Y(_1800_), .A(regs_14__30_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf3), );
  AOI21X1 AOI21X1_95 (.Y(_183_), .A(_1061__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf2), .C(_1800_), );
  NOR2X1 NOR2X1_104 (.Y(_1801_), .A(regs_14__31_), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf1), );
  AOI21X1 AOI21X1_96 (.Y(_184_), .A(_1063__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1769__bF_buf0), .C(_1801_), );
  INVX2 INVX2_161 (.Y(_1802_), .A(regs_13__0_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_105 (.Y(_1803_), .A(_1704__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1070__bF_buf8), );
  NAND2X1 NAND2X1_163 (.Y(_1804_), .A(wdata[0]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf7), );
  OAI21X1 OAI21X1_345 (.Y(_128_), .A(_1802_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf6), .C(_1804_), );
  INVX2 INVX2_162 (.Y(_1805_), .A(regs_13__1_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_164 (.Y(_1806_), .A(wdata[1]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf5), );
  OAI21X1 OAI21X1_346 (.Y(_139_), .A(_1805_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf4), .C(_1806_), );
  INVX2 INVX2_163 (.Y(_1807_), .A(regs_13__2_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_165 (.Y(_1808_), .A(wdata[2]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf3), );
  OAI21X1 OAI21X1_347 (.Y(_150_), .A(_1807_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf2), .C(_1808_), );
  INVX2 INVX2_164 (.Y(_1809_), .A(regs_13__3_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_166 (.Y(_1810_), .A(wdata[3]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf1), );
  OAI21X1 OAI21X1_348 (.Y(_153_), .A(_1809_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf0), .C(_1810_), );
  INVX2 INVX2_165 (.Y(_1811_), .A(regs_13__4_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_167 (.Y(_1812_), .A(wdata[4]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf7), );
  OAI21X1 OAI21X1_349 (.Y(_154_), .A(_1811_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf6), .C(_1812_), );
  INVX2 INVX2_166 (.Y(_1813_), .A(regs_13__5_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_168 (.Y(_1814_), .A(wdata[5]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf5), );
  OAI21X1 OAI21X1_350 (.Y(_155_), .A(_1813_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf4), .C(_1814_), );
  INVX2 INVX2_167 (.Y(_1815_), .A(regs_13__6_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_169 (.Y(_1816_), .A(wdata[6]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf3), );
  OAI21X1 OAI21X1_351 (.Y(_156_), .A(_1815_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf2), .C(_1816_), );
  INVX2 INVX2_168 (.Y(_1817_), .A(regs_13__7_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_170 (.Y(_1818_), .A(wdata[7]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf1), );
  OAI21X1 OAI21X1_352 (.Y(_157_), .A(_1817_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf0), .C(_1818_), );
  INVX2 INVX2_169 (.Y(_1819_), .A(regs_13__8_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_171 (.Y(_1820_), .A(wdata[8]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf7), );
  OAI21X1 OAI21X1_353 (.Y(_158_), .A(_1819_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf6), .C(_1820_), );
  INVX2 INVX2_170 (.Y(_1821_), .A(regs_13__9_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_172 (.Y(_1822_), .A(wdata[9]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf5), );
  OAI21X1 OAI21X1_354 (.Y(_159_), .A(_1821_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf4), .C(_1822_), );
  INVX2 INVX2_171 (.Y(_1823_), .A(regs_13__10_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_173 (.Y(_1824_), .A(wdata[10]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf3), );
  OAI21X1 OAI21X1_355 (.Y(_129_), .A(_1823_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf2), .C(_1824_), );
  INVX2 INVX2_172 (.Y(_1825_), .A(regs_13__11_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_174 (.Y(_1826_), .A(wdata[11]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf1), );
  OAI21X1 OAI21X1_356 (.Y(_130_), .A(_1825_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf0), .C(_1826_), );
  INVX2 INVX2_173 (.Y(_1827_), .A(regs_13__12_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_175 (.Y(_1828_), .A(wdata[12]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf7), );
  OAI21X1 OAI21X1_357 (.Y(_131_), .A(_1827_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf6), .C(_1828_), );
  INVX2 INVX2_174 (.Y(_1829_), .A(regs_13__13_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_176 (.Y(_1830_), .A(wdata[13]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf5), );
  OAI21X1 OAI21X1_358 (.Y(_132_), .A(_1829_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf4), .C(_1830_), );
  INVX2 INVX2_175 (.Y(_1831_), .A(regs_13__14_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_177 (.Y(_1832_), .A(wdata[14]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf3), );
  OAI21X1 OAI21X1_359 (.Y(_133_), .A(_1831_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf2), .C(_1832_), );
  INVX2 INVX2_176 (.Y(_1833_), .A(regs_13__15_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_178 (.Y(_1834_), .A(wdata[15]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf1), );
  OAI21X1 OAI21X1_360 (.Y(_134_), .A(_1833_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf0), .C(_1834_), );
  INVX2 INVX2_177 (.Y(_1835_), .A(regs_13__16_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_179 (.Y(_1836_), .A(wdata[16]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf7), );
  OAI21X1 OAI21X1_361 (.Y(_135_), .A(_1835_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf6), .C(_1836_), );
  INVX2 INVX2_178 (.Y(_1837_), .A(regs_13__17_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_180 (.Y(_1838_), .A(wdata[17]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf5), );
  OAI21X1 OAI21X1_362 (.Y(_136_), .A(_1837_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf4), .C(_1838_), );
  INVX2 INVX2_179 (.Y(_1839_), .A(regs_13__18_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_181 (.Y(_1840_), .A(wdata[18]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf3), );
  OAI21X1 OAI21X1_363 (.Y(_137_), .A(_1839_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf2), .C(_1840_), );
  INVX2 INVX2_180 (.Y(_1841_), .A(regs_13__19_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_182 (.Y(_1842_), .A(wdata[19]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf1), );
  OAI21X1 OAI21X1_364 (.Y(_138_), .A(_1841_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf0), .C(_1842_), );
  INVX2 INVX2_181 (.Y(_1843_), .A(regs_13__20_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_183 (.Y(_1844_), .A(wdata[20]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf7), );
  OAI21X1 OAI21X1_365 (.Y(_140_), .A(_1843_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf6), .C(_1844_), );
  INVX2 INVX2_182 (.Y(_1845_), .A(regs_13__21_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_184 (.Y(_1846_), .A(wdata[21]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf5), );
  OAI21X1 OAI21X1_366 (.Y(_141_), .A(_1845_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf4), .C(_1846_), );
  INVX2 INVX2_183 (.Y(_1847_), .A(regs_13__22_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_185 (.Y(_1848_), .A(wdata[22]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf3), );
  OAI21X1 OAI21X1_367 (.Y(_142_), .A(_1847_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf2), .C(_1848_), );
  INVX2 INVX2_184 (.Y(_1849_), .A(regs_13__23_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_186 (.Y(_1850_), .A(wdata[23]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf1), );
  OAI21X1 OAI21X1_368 (.Y(_143_), .A(_1849_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf0), .C(_1850_), );
  INVX2 INVX2_185 (.Y(_1851_), .A(regs_13__24_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_187 (.Y(_1852_), .A(wdata[24]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf7), );
  OAI21X1 OAI21X1_369 (.Y(_144_), .A(_1851_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf6), .C(_1852_), );
  INVX2 INVX2_186 (.Y(_1853_), .A(regs_13__25_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_188 (.Y(_1854_), .A(wdata[25]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf5), );
  OAI21X1 OAI21X1_370 (.Y(_145_), .A(_1853_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf4), .C(_1854_), );
  INVX2 INVX2_187 (.Y(_1855_), .A(regs_13__26_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_189 (.Y(_1856_), .A(wdata[26]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf3), );
  OAI21X1 OAI21X1_371 (.Y(_146_), .A(_1855_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf2), .C(_1856_), );
  INVX2 INVX2_188 (.Y(_1857_), .A(regs_13__27_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_190 (.Y(_1858_), .A(wdata[27]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf1), );
  OAI21X1 OAI21X1_372 (.Y(_147_), .A(_1857_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf0), .C(_1858_), );
  INVX2 INVX2_189 (.Y(_1859_), .A(regs_13__28_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_191 (.Y(_1860_), .A(wdata[28]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf7), );
  OAI21X1 OAI21X1_373 (.Y(_148_), .A(_1859_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf6), .C(_1860_), );
  INVX2 INVX2_190 (.Y(_1861_), .A(regs_13__29_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_192 (.Y(_1862_), .A(wdata[29]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf5), );
  OAI21X1 OAI21X1_374 (.Y(_149_), .A(_1861_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf4), .C(_1862_), );
  INVX2 INVX2_191 (.Y(_1863_), .A(regs_13__30_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_193 (.Y(_1864_), .A(wdata[30]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf3), );
  OAI21X1 OAI21X1_375 (.Y(_151_), .A(_1863_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf2), .C(_1864_), );
  INVX2 INVX2_192 (.Y(_1865_), .A(regs_13__31_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_194 (.Y(_1866_), .A(wdata[31]), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf1), );
  OAI21X1 OAI21X1_376 (.Y(_152_), .A(_1865_), .gnd(gnd), .vdd(vdd), .B(_1803__bF_buf0), .C(_1866_), );
  OR2X2 OR2X2_6 (.Y(_1867_), .A(_1704__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf10), );
  OAI21X1 OAI21X1_377 (.Y(_1868_), .A(_1704__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf9), .C(regs_12__0_), );
  OAI21X1 OAI21X1_378 (.Y(_96_), .A(_1867__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_992__bF_buf2), .C(_1868_), );
  OAI21X1 OAI21X1_379 (.Y(_1869_), .A(_1704__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf8), .C(regs_12__1_), );
  OAI21X1 OAI21X1_380 (.Y(_107_), .A(_1867__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1003__bF_buf2), .C(_1869_), );
  OAI21X1 OAI21X1_381 (.Y(_1870_), .A(_1704__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf7), .C(regs_12__2_), );
  OAI21X1 OAI21X1_382 (.Y(_118_), .A(_1867__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1005__bF_buf2), .C(_1870_), );
  OAI21X1 OAI21X1_383 (.Y(_1871_), .A(_1704__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf6), .C(regs_12__3_), );
  OAI21X1 OAI21X1_384 (.Y(_121_), .A(_1867__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1007__bF_buf2), .C(_1871_), );
  OAI21X1 OAI21X1_385 (.Y(_1872_), .A(_1704__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf5), .C(regs_12__4_), );
  OAI21X1 OAI21X1_386 (.Y(_122_), .A(_1867__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1009__bF_buf1), .C(_1872_), );
  OAI21X1 OAI21X1_387 (.Y(_1873_), .A(_1704__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf4), .C(regs_12__5_), );
  OAI21X1 OAI21X1_388 (.Y(_123_), .A(_1867__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1011__bF_buf1), .C(_1873_), );
  OAI21X1 OAI21X1_389 (.Y(_1874_), .A(_1704__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf3), .C(regs_12__6_), );
  OAI21X1 OAI21X1_390 (.Y(_124_), .A(_1867__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1013__bF_buf1), .C(_1874_), );
  OAI21X1 OAI21X1_391 (.Y(_1875_), .A(_1704__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf2), .C(regs_12__7_), );
  OAI21X1 OAI21X1_392 (.Y(_125_), .A(_1867__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1015__bF_buf1), .C(_1875_), );
  OAI21X1 OAI21X1_393 (.Y(_1876_), .A(_1704__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf1), .C(regs_12__8_), );
  OAI21X1 OAI21X1_394 (.Y(_126_), .A(_1867__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1017__bF_buf1), .C(_1876_), );
  OAI21X1 OAI21X1_395 (.Y(_1877_), .A(_1704__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf0), .C(regs_12__9_), );
  OAI21X1 OAI21X1_396 (.Y(_127_), .A(_1867__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1019__bF_buf1), .C(_1877_), );
  OAI21X1 OAI21X1_397 (.Y(_1878_), .A(_1704__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf14), .C(regs_12__10_), );
  OAI21X1 OAI21X1_398 (.Y(_97_), .A(_1867__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1021__bF_buf1), .C(_1878_), );
  OAI21X1 OAI21X1_399 (.Y(_1879_), .A(_1704__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf13), .C(regs_12__11_), );
  OAI21X1 OAI21X1_400 (.Y(_98_), .A(_1867__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1023__bF_buf1), .C(_1879_), );
  OAI21X1 OAI21X1_401 (.Y(_1880_), .A(_1704__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf12), .C(regs_12__12_), );
  OAI21X1 OAI21X1_402 (.Y(_99_), .A(_1867__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1025__bF_buf1), .C(_1880_), );
  OAI21X1 OAI21X1_403 (.Y(_1881_), .A(_1704__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf11), .C(regs_12__13_), );
  OAI21X1 OAI21X1_404 (.Y(_100_), .A(_1867__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1027__bF_buf1), .C(_1881_), );
  OAI21X1 OAI21X1_405 (.Y(_1882_), .A(_1704__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf10), .C(regs_12__14_), );
  OAI21X1 OAI21X1_406 (.Y(_101_), .A(_1867__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1029__bF_buf1), .C(_1882_), );
  OAI21X1 OAI21X1_407 (.Y(_1883_), .A(_1704__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf9), .C(regs_12__15_), );
  OAI21X1 OAI21X1_408 (.Y(_102_), .A(_1867__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1031__bF_buf1), .C(_1883_), );
  OAI21X1 OAI21X1_409 (.Y(_1884_), .A(_1704__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf8), .C(regs_12__16_), );
  OAI21X1 OAI21X1_410 (.Y(_103_), .A(_1867__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1033__bF_buf1), .C(_1884_), );
  OAI21X1 OAI21X1_411 (.Y(_1885_), .A(_1704__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf7), .C(regs_12__17_), );
  OAI21X1 OAI21X1_412 (.Y(_104_), .A(_1867__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1035__bF_buf1), .C(_1885_), );
  OAI21X1 OAI21X1_413 (.Y(_1886_), .A(_1704__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf6), .C(regs_12__18_), );
  OAI21X1 OAI21X1_414 (.Y(_105_), .A(_1867__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1037__bF_buf1), .C(_1886_), );
  OAI21X1 OAI21X1_415 (.Y(_1887_), .A(_1704__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf5), .C(regs_12__19_), );
  OAI21X1 OAI21X1_416 (.Y(_106_), .A(_1867__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1039__bF_buf1), .C(_1887_), );
  OAI21X1 OAI21X1_417 (.Y(_1888_), .A(_1704__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf4), .C(regs_12__20_), );
  OAI21X1 OAI21X1_418 (.Y(_108_), .A(_1867__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1041__bF_buf1), .C(_1888_), );
  OAI21X1 OAI21X1_419 (.Y(_1889_), .A(_1704__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf3), .C(regs_12__21_), );
  OAI21X1 OAI21X1_420 (.Y(_109_), .A(_1867__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1043__bF_buf1), .C(_1889_), );
  OAI21X1 OAI21X1_421 (.Y(_1890_), .A(_1704__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf2), .C(regs_12__22_), );
  OAI21X1 OAI21X1_422 (.Y(_110_), .A(_1867__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1045__bF_buf1), .C(_1890_), );
  OAI21X1 OAI21X1_423 (.Y(_1891_), .A(_1704__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf1), .C(regs_12__23_), );
  OAI21X1 OAI21X1_424 (.Y(_111_), .A(_1867__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1047__bF_buf1), .C(_1891_), );
  OAI21X1 OAI21X1_425 (.Y(_1892_), .A(_1704__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf0), .C(regs_12__24_), );
  OAI21X1 OAI21X1_426 (.Y(_112_), .A(_1867__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1049__bF_buf1), .C(_1892_), );
  OAI21X1 OAI21X1_427 (.Y(_1893_), .A(_1704__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf14), .C(regs_12__25_), );
  OAI21X1 OAI21X1_428 (.Y(_113_), .A(_1867__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1051__bF_buf1), .C(_1893_), );
  OAI21X1 OAI21X1_429 (.Y(_1894_), .A(_1704__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf13), .C(regs_12__26_), );
  OAI21X1 OAI21X1_430 (.Y(_114_), .A(_1867__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1053__bF_buf1), .C(_1894_), );
  OAI21X1 OAI21X1_431 (.Y(_1895_), .A(_1704__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf12), .C(regs_12__27_), );
  OAI21X1 OAI21X1_432 (.Y(_115_), .A(_1867__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1055__bF_buf1), .C(_1895_), );
  OAI21X1 OAI21X1_433 (.Y(_1896_), .A(_1704__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf11), .C(regs_12__28_), );
  OAI21X1 OAI21X1_434 (.Y(_116_), .A(_1867__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1057__bF_buf1), .C(_1896_), );
  OAI21X1 OAI21X1_435 (.Y(_1897_), .A(_1704__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf10), .C(regs_12__29_), );
  OAI21X1 OAI21X1_436 (.Y(_117_), .A(_1867__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1059__bF_buf1), .C(_1897_), );
  OAI21X1 OAI21X1_437 (.Y(_1898_), .A(_1704__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf9), .C(regs_12__30_), );
  OAI21X1 OAI21X1_438 (.Y(_119_), .A(_1867__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1061__bF_buf1), .C(_1898_), );
  OAI21X1 OAI21X1_439 (.Y(_1899_), .A(_1704__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf8), .C(regs_12__31_), );
  OAI21X1 OAI21X1_440 (.Y(_120_), .A(_1867__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1063__bF_buf1), .C(_1899_), );
  INVX2 INVX2_193 (.Y(_1900_), .A(regs_11__0_), .gnd(gnd), .vdd(vdd), );
  OR2X2 OR2X2_7 (.Y(_1901_), .A(_1703_), .gnd(gnd), .vdd(vdd), .B(_1139_), );
  NOR2X1 NOR2X1_106 (.Y(_1902_), .A(_1142__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1901__bF_buf5), );
  NAND2X1 NAND2X1_195 (.Y(_1903_), .A(wdata[0]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf7), );
  OAI21X1 OAI21X1_441 (.Y(_64_), .A(_1900_), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf6), .C(_1903_), );
  INVX2 INVX2_194 (.Y(_1904_), .A(regs_11__1_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_196 (.Y(_1905_), .A(wdata[1]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf5), );
  OAI21X1 OAI21X1_442 (.Y(_75_), .A(_1904_), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf4), .C(_1905_), );
  INVX2 INVX2_195 (.Y(_1906_), .A(regs_11__2_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_197 (.Y(_1907_), .A(wdata[2]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf3), );
  OAI21X1 OAI21X1_443 (.Y(_86_), .A(_1906_), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf2), .C(_1907_), );
  INVX2 INVX2_196 (.Y(_1908_), .A(regs_11__3_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_198 (.Y(_1909_), .A(wdata[3]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf1), );
  OAI21X1 OAI21X1_444 (.Y(_89_), .A(_1908_), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf0), .C(_1909_), );
  INVX2 INVX2_197 (.Y(_1910_), .A(regs_11__4_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_199 (.Y(_1911_), .A(wdata[4]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf7), );
  OAI21X1 OAI21X1_445 (.Y(_90_), .A(_1910_), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf6), .C(_1911_), );
  INVX2 INVX2_198 (.Y(_1912_), .A(regs_11__5_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_200 (.Y(_1913_), .A(wdata[5]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf5), );
  OAI21X1 OAI21X1_446 (.Y(_91_), .A(_1912_), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf4), .C(_1913_), );
  INVX2 INVX2_199 (.Y(_1914_), .A(regs_11__6_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_201 (.Y(_1915_), .A(wdata[6]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf3), );
  OAI21X1 OAI21X1_447 (.Y(_92_), .A(_1914_), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf2), .C(_1915_), );
  INVX2 INVX2_200 (.Y(_1916_), .A(regs_11__7_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_202 (.Y(_1917_), .A(wdata[7]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf1), );
  OAI21X1 OAI21X1_448 (.Y(_93_), .A(_1916_), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf0), .C(_1917_), );
  INVX2 INVX2_201 (.Y(_1918_), .A(regs_11__8_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_203 (.Y(_1919_), .A(wdata[8]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf7), );
  OAI21X1 OAI21X1_449 (.Y(_94_), .A(_1918_), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf6), .C(_1919_), );
  INVX2 INVX2_202 (.Y(_1920_), .A(regs_11__9_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_204 (.Y(_1921_), .A(wdata[9]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf5), );
  OAI21X1 OAI21X1_450 (.Y(_95_), .A(_1920_), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf4), .C(_1921_), );
  INVX2 INVX2_203 (.Y(_1922_), .A(regs_11__10_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_205 (.Y(_1923_), .A(wdata[10]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf3), );
  OAI21X1 OAI21X1_451 (.Y(_65_), .A(_1922_), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf2), .C(_1923_), );
  INVX2 INVX2_204 (.Y(_1924_), .A(regs_11__11_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_206 (.Y(_1925_), .A(wdata[11]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf1), );
  OAI21X1 OAI21X1_452 (.Y(_66_), .A(_1924_), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf0), .C(_1925_), );
  INVX2 INVX2_205 (.Y(_1926_), .A(regs_11__12_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_207 (.Y(_1927_), .A(wdata[12]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf7), );
  OAI21X1 OAI21X1_453 (.Y(_67_), .A(_1926_), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf6), .C(_1927_), );
  INVX2 INVX2_206 (.Y(_1928_), .A(regs_11__13_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_208 (.Y(_1929_), .A(wdata[13]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf5), );
  OAI21X1 OAI21X1_454 (.Y(_68_), .A(_1928_), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf4), .C(_1929_), );
  INVX2 INVX2_207 (.Y(_1930_), .A(regs_11__14_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_209 (.Y(_1931_), .A(wdata[14]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf3), );
  OAI21X1 OAI21X1_455 (.Y(_69_), .A(_1930_), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf2), .C(_1931_), );
  INVX2 INVX2_208 (.Y(_1932_), .A(regs_11__15_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_210 (.Y(_1933_), .A(wdata[15]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf1), );
  OAI21X1 OAI21X1_456 (.Y(_70_), .A(_1932_), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf0), .C(_1933_), );
  INVX2 INVX2_209 (.Y(_1934_), .A(regs_11__16_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_211 (.Y(_1935_), .A(wdata[16]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf7), );
  OAI21X1 OAI21X1_457 (.Y(_71_), .A(_1934_), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf6), .C(_1935_), );
  INVX2 INVX2_210 (.Y(_1936_), .A(regs_11__17_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_212 (.Y(_1937_), .A(wdata[17]), .gnd(gnd), .vdd(vdd), .B(_1902__bF_buf5), );
  BUFX2 BUFX2_1 (.Y(rdata1[0]), .A(_5511__0_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_2 (.Y(rdata1[1]), .A(_5511__1_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_3 (.Y(rdata1[2]), .A(_5511__2_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_4 (.Y(rdata1[3]), .A(_5511__3_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_5 (.Y(rdata1[4]), .A(_5511__4_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_6 (.Y(rdata1[5]), .A(_5511__5_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_7 (.Y(rdata1[6]), .A(_5511__6_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_8 (.Y(rdata1[7]), .A(_5511__7_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_9 (.Y(rdata1[8]), .A(_5511__8_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_10 (.Y(rdata1[9]), .A(_5511__9_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_11 (.Y(rdata1[10]), .A(_5511__10_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_12 (.Y(rdata1[11]), .A(_5511__11_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_13 (.Y(rdata1[12]), .A(_5511__12_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_14 (.Y(rdata1[13]), .A(_5511__13_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_15 (.Y(rdata1[14]), .A(_5511__14_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_16 (.Y(rdata1[15]), .A(_5511__15_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_17 (.Y(rdata1[16]), .A(_5511__16_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_18 (.Y(rdata1[17]), .A(_5511__17_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_19 (.Y(rdata1[18]), .A(_5511__18_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_20 (.Y(rdata1[19]), .A(_5511__19_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_21 (.Y(rdata1[20]), .A(_5511__20_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_22 (.Y(rdata1[21]), .A(_5511__21_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_23 (.Y(rdata1[22]), .A(_5511__22_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_24 (.Y(rdata1[23]), .A(_5511__23_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_25 (.Y(rdata1[24]), .A(_5511__24_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_26 (.Y(rdata1[25]), .A(_5511__25_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_27 (.Y(rdata1[26]), .A(_5511__26_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_28 (.Y(rdata1[27]), .A(_5511__27_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_29 (.Y(rdata1[28]), .A(_5511__28_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_30 (.Y(rdata1[29]), .A(_5511__29_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_31 (.Y(rdata1[30]), .A(_5511__30_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_32 (.Y(rdata1[31]), .A(_5511__31_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_33 (.Y(rdata2[0]), .A(_5512__0_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_34 (.Y(rdata2[1]), .A(_5512__1_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_35 (.Y(rdata2[2]), .A(_5512__2_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_36 (.Y(rdata2[3]), .A(_5512__3_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_37 (.Y(rdata2[4]), .A(_5512__4_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_38 (.Y(rdata2[5]), .A(_5512__5_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_39 (.Y(rdata2[6]), .A(_5512__6_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_40 (.Y(rdata2[7]), .A(_5512__7_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_41 (.Y(rdata2[8]), .A(_5512__8_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_42 (.Y(rdata2[9]), .A(_5512__9_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_43 (.Y(rdata2[10]), .A(_5512__10_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_44 (.Y(rdata2[11]), .A(_5512__11_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_45 (.Y(rdata2[12]), .A(_5512__12_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_46 (.Y(rdata2[13]), .A(_5512__13_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_47 (.Y(rdata2[14]), .A(_5512__14_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_48 (.Y(rdata2[15]), .A(_5512__15_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_49 (.Y(rdata2[16]), .A(_5512__16_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_50 (.Y(rdata2[17]), .A(_5512__17_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_51 (.Y(rdata2[18]), .A(_5512__18_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_52 (.Y(rdata2[19]), .A(_5512__19_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_53 (.Y(rdata2[20]), .A(_5512__20_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_54 (.Y(rdata2[21]), .A(_5512__21_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_55 (.Y(rdata2[22]), .A(_5512__22_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_56 (.Y(rdata2[23]), .A(_5512__23_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_57 (.Y(rdata2[24]), .A(_5512__24_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_58 (.Y(rdata2[25]), .A(_5512__25_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_59 (.Y(rdata2[26]), .A(_5512__26_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_60 (.Y(rdata2[27]), .A(_5512__27_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_61 (.Y(rdata2[28]), .A(_5512__28_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_62 (.Y(rdata2[29]), .A(_5512__29_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_63 (.Y(rdata2[30]), .A(_5512__30_), .gnd(gnd), .vdd(vdd), );
  BUFX2 BUFX2_64 (.Y(rdata2[31]), .A(_5512__31_), .gnd(gnd), .vdd(vdd), );
  DFFPOSX1 DFFPOSX1_1 (.Q(regs_1__0_), .gnd(gnd), .vdd(vdd), .D(_352_), .CLK(clock_bf2__0), );
  DFFPOSX1 DFFPOSX1_2 (.Q(regs_1__1_), .gnd(gnd), .vdd(vdd), .D(_363_), .CLK(clock_bf2__11), );
  DFFPOSX1 DFFPOSX1_3 (.Q(regs_1__2_), .gnd(gnd), .vdd(vdd), .D(_374_), .CLK(random_clk_bf3__401), );
  DFFPOSX1 DFFPOSX1_4 (.Q(regs_1__3_), .gnd(gnd), .vdd(vdd), .D(_377_), .CLK(random_clk_bf3__621), );
  DFFPOSX1 DFFPOSX1_5 (.Q(regs_1__4_), .gnd(gnd), .vdd(vdd), .D(_378_), .CLK(random_clk_bf3__841), );
  DFFPOSX1 DFFPOSX1_6 (.Q(regs_1__5_), .gnd(gnd), .vdd(vdd), .D(_379_), .CLK(random_clk_bf3__1061), );
  DFFPOSX1 DFFPOSX1_7 (.Q(regs_1__6_), .gnd(gnd), .vdd(vdd), .D(_380_), .CLK(random_clk_bf3__1281), );
  DFFPOSX1 DFFPOSX1_8 (.Q(regs_1__7_), .gnd(gnd), .vdd(vdd), .D(_381_), .CLK(random_clk_bf3__1501), );
  DFFPOSX1 DFFPOSX1_9 (.Q(regs_1__8_), .gnd(gnd), .vdd(vdd), .D(_382_), .CLK(random_clk_bf3__1721), );
  DFFPOSX1 DFFPOSX1_10 (.Q(regs_1__9_), .gnd(gnd), .vdd(vdd), .D(_383_), .CLK(random_clk_bf3__1), );
  DFFPOSX1 DFFPOSX1_11 (.Q(regs_1__10_), .gnd(gnd), .vdd(vdd), .D(_353_), .CLK(random_clk_bf3__201), );
  DFFPOSX1 DFFPOSX1_12 (.Q(regs_1__11_), .gnd(gnd), .vdd(vdd), .D(_354_), .CLK(random_clk_bf3__421), );
  DFFPOSX1 DFFPOSX1_13 (.Q(regs_1__12_), .gnd(gnd), .vdd(vdd), .D(_355_), .CLK(random_clk_bf3__641), );
  DFFPOSX1 DFFPOSX1_14 (.Q(regs_1__13_), .gnd(gnd), .vdd(vdd), .D(_356_), .CLK(random_clk_bf3__861), );
  DFFPOSX1 DFFPOSX1_15 (.Q(regs_1__14_), .gnd(gnd), .vdd(vdd), .D(_357_), .CLK(random_clk_bf3__1081), );
  DFFPOSX1 DFFPOSX1_16 (.Q(regs_1__15_), .gnd(gnd), .vdd(vdd), .D(_358_), .CLK(random_clk_bf3__1301), );
  DFFPOSX1 DFFPOSX1_17 (.Q(regs_1__16_), .gnd(gnd), .vdd(vdd), .D(_359_), .CLK(random_clk_bf3__1521), );
  DFFPOSX1 DFFPOSX1_18 (.Q(regs_1__17_), .gnd(gnd), .vdd(vdd), .D(_360_), .CLK(random_clk_bf3__1741), );
  DFFPOSX1 DFFPOSX1_19 (.Q(regs_1__18_), .gnd(gnd), .vdd(vdd), .D(_361_), .CLK(random_clk_bf3__21), );
  DFFPOSX1 DFFPOSX1_20 (.Q(regs_1__19_), .gnd(gnd), .vdd(vdd), .D(_362_), .CLK(random_clk_bf3__221), );
  DFFPOSX1 DFFPOSX1_21 (.Q(regs_1__20_), .gnd(gnd), .vdd(vdd), .D(_364_), .CLK(random_clk_bf3__441), );
  DFFPOSX1 DFFPOSX1_22 (.Q(regs_1__21_), .gnd(gnd), .vdd(vdd), .D(_365_), .CLK(random_clk_bf3__661), );
  DFFPOSX1 DFFPOSX1_23 (.Q(regs_1__22_), .gnd(gnd), .vdd(vdd), .D(_366_), .CLK(random_clk_bf3__881), );
  DFFPOSX1 DFFPOSX1_24 (.Q(regs_1__23_), .gnd(gnd), .vdd(vdd), .D(_367_), .CLK(random_clk_bf3__1101), );
  DFFPOSX1 DFFPOSX1_25 (.Q(regs_1__24_), .gnd(gnd), .vdd(vdd), .D(_368_), .CLK(random_clk_bf3__1321), );
  DFFPOSX1 DFFPOSX1_26 (.Q(regs_1__25_), .gnd(gnd), .vdd(vdd), .D(_369_), .CLK(random_clk_bf3__1541), );
  DFFPOSX1 DFFPOSX1_27 (.Q(regs_1__26_), .gnd(gnd), .vdd(vdd), .D(_370_), .CLK(random_clk_bf3__1761), );
  DFFPOSX1 DFFPOSX1_28 (.Q(regs_1__27_), .gnd(gnd), .vdd(vdd), .D(_371_), .CLK(random_clk_bf3__41), );
  DFFPOSX1 DFFPOSX1_29 (.Q(regs_1__28_), .gnd(gnd), .vdd(vdd), .D(_372_), .CLK(random_clk_bf3__241), );
  DFFPOSX1 DFFPOSX1_30 (.Q(regs_1__29_), .gnd(gnd), .vdd(vdd), .D(_373_), .CLK(random_clk_bf3__461), );
  DFFPOSX1 DFFPOSX1_31 (.Q(regs_1__30_), .gnd(gnd), .vdd(vdd), .D(_375_), .CLK(random_clk_bf3__681), );
  DFFPOSX1 DFFPOSX1_32 (.Q(regs_1__31_), .gnd(gnd), .vdd(vdd), .D(_376_), .CLK(random_clk_bf3__901), );
  DFFPOSX1 DFFPOSX1_33 (.Q(regs_0__0_), .gnd(gnd), .vdd(vdd), .D(_0_), .CLK(random_clk_bf3__1121), );
  DFFPOSX1 DFFPOSX1_34 (.Q(regs_0__1_), .gnd(gnd), .vdd(vdd), .D(_11_), .CLK(random_clk_bf3__1341), );
  DFFPOSX1 DFFPOSX1_35 (.Q(regs_0__2_), .gnd(gnd), .vdd(vdd), .D(_22_), .CLK(random_clk_bf3__1561), );
  DFFPOSX1 DFFPOSX1_36 (.Q(regs_0__3_), .gnd(gnd), .vdd(vdd), .D(_25_), .CLK(random_clk_bf3__1781), );
  DFFPOSX1 DFFPOSX1_37 (.Q(regs_0__4_), .gnd(gnd), .vdd(vdd), .D(_26_), .CLK(random_clk_bf3__61), );
  DFFPOSX1 DFFPOSX1_38 (.Q(regs_0__5_), .gnd(gnd), .vdd(vdd), .D(_27_), .CLK(random_clk_bf3__261), );
  DFFPOSX1 DFFPOSX1_39 (.Q(regs_0__6_), .gnd(gnd), .vdd(vdd), .D(_28_), .CLK(random_clk_bf3__481), );
  DFFPOSX1 DFFPOSX1_40 (.Q(regs_0__7_), .gnd(gnd), .vdd(vdd), .D(_29_), .CLK(random_clk_bf3__701), );
  DFFPOSX1 DFFPOSX1_41 (.Q(regs_0__8_), .gnd(gnd), .vdd(vdd), .D(_30_), .CLK(random_clk_bf3__921), );
  DFFPOSX1 DFFPOSX1_42 (.Q(regs_0__9_), .gnd(gnd), .vdd(vdd), .D(_31_), .CLK(random_clk_bf3__1141), );
  DFFPOSX1 DFFPOSX1_43 (.Q(regs_0__10_), .gnd(gnd), .vdd(vdd), .D(_1_), .CLK(random_clk_bf3__1361), );
  DFFPOSX1 DFFPOSX1_44 (.Q(regs_0__11_), .gnd(gnd), .vdd(vdd), .D(_2_), .CLK(random_clk_bf3__1581), );
  DFFPOSX1 DFFPOSX1_45 (.Q(regs_0__12_), .gnd(gnd), .vdd(vdd), .D(_3_), .CLK(random_clk_bf3__1801), );
  DFFPOSX1 DFFPOSX1_46 (.Q(regs_0__13_), .gnd(gnd), .vdd(vdd), .D(_4_), .CLK(random_clk_bf3__81), );
  DFFPOSX1 DFFPOSX1_47 (.Q(regs_0__14_), .gnd(gnd), .vdd(vdd), .D(_5_), .CLK(random_clk_bf3__281), );
  DFFPOSX1 DFFPOSX1_48 (.Q(regs_0__15_), .gnd(gnd), .vdd(vdd), .D(_6_), .CLK(random_clk_bf3__501), );
  DFFPOSX1 DFFPOSX1_49 (.Q(regs_0__16_), .gnd(gnd), .vdd(vdd), .D(_7_), .CLK(random_clk_bf3__721), );
  DFFPOSX1 DFFPOSX1_50 (.Q(regs_0__17_), .gnd(gnd), .vdd(vdd), .D(_8_), .CLK(random_clk_bf3__941), );
  DFFPOSX1 DFFPOSX1_51 (.Q(regs_0__18_), .gnd(gnd), .vdd(vdd), .D(_9_), .CLK(random_clk_bf3__1161), );
  DFFPOSX1 DFFPOSX1_52 (.Q(regs_0__19_), .gnd(gnd), .vdd(vdd), .D(_10_), .CLK(random_clk_bf3__1381), );
  DFFPOSX1 DFFPOSX1_53 (.Q(regs_0__20_), .gnd(gnd), .vdd(vdd), .D(_12_), .CLK(random_clk_bf3__1601), );
  DFFPOSX1 DFFPOSX1_54 (.Q(regs_0__21_), .gnd(gnd), .vdd(vdd), .D(_13_), .CLK(random_clk_bf3__1821), );
  DFFPOSX1 DFFPOSX1_55 (.Q(regs_0__22_), .gnd(gnd), .vdd(vdd), .D(_14_), .CLK(random_clk_bf3__101), );
  DFFPOSX1 DFFPOSX1_56 (.Q(regs_0__23_), .gnd(gnd), .vdd(vdd), .D(_15_), .CLK(random_clk_bf3__301), );
  DFFPOSX1 DFFPOSX1_57 (.Q(regs_0__24_), .gnd(gnd), .vdd(vdd), .D(_16_), .CLK(random_clk_bf3__521), );
  DFFPOSX1 DFFPOSX1_58 (.Q(regs_0__25_), .gnd(gnd), .vdd(vdd), .D(_17_), .CLK(random_clk_bf3__741), );
  DFFPOSX1 DFFPOSX1_59 (.Q(regs_0__26_), .gnd(gnd), .vdd(vdd), .D(_18_), .CLK(random_clk_bf3__961), );
  DFFPOSX1 DFFPOSX1_60 (.Q(regs_0__27_), .gnd(gnd), .vdd(vdd), .D(_19_), .CLK(random_clk_bf3__1181), );
  DFFPOSX1 DFFPOSX1_61 (.Q(regs_0__28_), .gnd(gnd), .vdd(vdd), .D(_20_), .CLK(random_clk_bf3__1401), );
  DFFPOSX1 DFFPOSX1_62 (.Q(regs_0__29_), .gnd(gnd), .vdd(vdd), .D(_21_), .CLK(random_clk_bf3__1621), );
  DFFPOSX1 DFFPOSX1_63 (.Q(regs_0__30_), .gnd(gnd), .vdd(vdd), .D(_23_), .CLK(random_clk_bf3__1841), );
  DFFPOSX1 DFFPOSX1_64 (.Q(regs_0__31_), .gnd(gnd), .vdd(vdd), .D(_24_), .CLK(random_clk_bf3__121), );
  DFFPOSX1 DFFPOSX1_65 (.Q(regs_28__0_), .gnd(gnd), .vdd(vdd), .D(_640_), .CLK(random_clk_bf3__321), );
  DFFPOSX1 DFFPOSX1_66 (.Q(regs_28__1_), .gnd(gnd), .vdd(vdd), .D(_651_), .CLK(random_clk_bf3__541), );
  DFFPOSX1 DFFPOSX1_67 (.Q(regs_28__2_), .gnd(gnd), .vdd(vdd), .D(_662_), .CLK(random_clk_bf3__761), );
  DFFPOSX1 DFFPOSX1_68 (.Q(regs_28__3_), .gnd(gnd), .vdd(vdd), .D(_665_), .CLK(random_clk_bf3__981), );
  DFFPOSX1 DFFPOSX1_69 (.Q(regs_28__4_), .gnd(gnd), .vdd(vdd), .D(_666_), .CLK(random_clk_bf3__1201), );
  DFFPOSX1 DFFPOSX1_70 (.Q(regs_28__5_), .gnd(gnd), .vdd(vdd), .D(_667_), .CLK(random_clk_bf3__1421), );
  DFFPOSX1 DFFPOSX1_71 (.Q(regs_28__6_), .gnd(gnd), .vdd(vdd), .D(_668_), .CLK(random_clk_bf3__1641), );
  DFFPOSX1 DFFPOSX1_72 (.Q(regs_28__7_), .gnd(gnd), .vdd(vdd), .D(_669_), .CLK(random_clk_bf3__1861), );
  DFFPOSX1 DFFPOSX1_73 (.Q(regs_28__8_), .gnd(gnd), .vdd(vdd), .D(_670_), .CLK(random_clk_bf3__141), );
  DFFPOSX1 DFFPOSX1_74 (.Q(regs_28__9_), .gnd(gnd), .vdd(vdd), .D(_671_), .CLK(random_clk_bf3__341), );
  DFFPOSX1 DFFPOSX1_75 (.Q(regs_28__10_), .gnd(gnd), .vdd(vdd), .D(_641_), .CLK(random_clk_bf3__561), );
  DFFPOSX1 DFFPOSX1_76 (.Q(regs_28__11_), .gnd(gnd), .vdd(vdd), .D(_642_), .CLK(random_clk_bf3__781), );
  DFFPOSX1 DFFPOSX1_77 (.Q(regs_28__12_), .gnd(gnd), .vdd(vdd), .D(_643_), .CLK(random_clk_bf3__1001), );
  DFFPOSX1 DFFPOSX1_78 (.Q(regs_28__13_), .gnd(gnd), .vdd(vdd), .D(_644_), .CLK(random_clk_bf3__1221), );
  DFFPOSX1 DFFPOSX1_79 (.Q(regs_28__14_), .gnd(gnd), .vdd(vdd), .D(_645_), .CLK(random_clk_bf3__1441), );
  DFFPOSX1 DFFPOSX1_80 (.Q(regs_28__15_), .gnd(gnd), .vdd(vdd), .D(_646_), .CLK(random_clk_bf3__1661), );
  DFFPOSX1 DFFPOSX1_81 (.Q(regs_28__16_), .gnd(gnd), .vdd(vdd), .D(_647_), .CLK(random_clk_bf3__1881), );
  DFFPOSX1 DFFPOSX1_82 (.Q(regs_28__17_), .gnd(gnd), .vdd(vdd), .D(_648_), .CLK(random_clk_bf3__161), );
  DFFPOSX1 DFFPOSX1_83 (.Q(regs_28__18_), .gnd(gnd), .vdd(vdd), .D(_649_), .CLK(random_clk_bf3__361), );
  DFFPOSX1 DFFPOSX1_84 (.Q(regs_28__19_), .gnd(gnd), .vdd(vdd), .D(_650_), .CLK(random_clk_bf3__581), );
  DFFPOSX1 DFFPOSX1_85 (.Q(regs_28__20_), .gnd(gnd), .vdd(vdd), .D(_652_), .CLK(random_clk_bf3__801), );
  DFFPOSX1 DFFPOSX1_86 (.Q(regs_28__21_), .gnd(gnd), .vdd(vdd), .D(_653_), .CLK(random_clk_bf3__1021), );
  DFFPOSX1 DFFPOSX1_87 (.Q(regs_28__22_), .gnd(gnd), .vdd(vdd), .D(_654_), .CLK(random_clk_bf3__1241), );
  DFFPOSX1 DFFPOSX1_88 (.Q(regs_28__23_), .gnd(gnd), .vdd(vdd), .D(_655_), .CLK(random_clk_bf3__1461), );
  DFFPOSX1 DFFPOSX1_89 (.Q(regs_28__24_), .gnd(gnd), .vdd(vdd), .D(_656_), .CLK(random_clk_bf3__1681), );
  DFFPOSX1 DFFPOSX1_90 (.Q(regs_28__25_), .gnd(gnd), .vdd(vdd), .D(_657_), .CLK(random_clk_bf3__1901), );
  DFFPOSX1 DFFPOSX1_91 (.Q(regs_28__26_), .gnd(gnd), .vdd(vdd), .D(_658_), .CLK(random_clk_bf3__181), );
  DFFPOSX1 DFFPOSX1_92 (.Q(regs_28__27_), .gnd(gnd), .vdd(vdd), .D(_659_), .CLK(random_clk_bf3__381), );
  DFFPOSX1 DFFPOSX1_93 (.Q(regs_28__28_), .gnd(gnd), .vdd(vdd), .D(_660_), .CLK(random_clk_bf3__601), );
  DFFPOSX1 DFFPOSX1_94 (.Q(regs_28__29_), .gnd(gnd), .vdd(vdd), .D(_661_), .CLK(random_clk_bf3__821), );
  DFFPOSX1 DFFPOSX1_95 (.Q(regs_28__30_), .gnd(gnd), .vdd(vdd), .D(_663_), .CLK(random_clk_bf3__1041), );
  DFFPOSX1 DFFPOSX1_96 (.Q(regs_28__31_), .gnd(gnd), .vdd(vdd), .D(_664_), .CLK(random_clk_bf3__1261), );
  DFFPOSX1 DFFPOSX1_97 (.Q(regs_30__0_), .gnd(gnd), .vdd(vdd), .D(_736_), .CLK(random_clk_bf3__1481), );
  DFFPOSX1 DFFPOSX1_98 (.Q(regs_30__1_), .gnd(gnd), .vdd(vdd), .D(_747_), .CLK(random_clk_bf3__1701), );
  DFFPOSX1 DFFPOSX1_99 (.Q(regs_30__2_), .gnd(gnd), .vdd(vdd), .D(_758_), .CLK(clock_bf2__22), );
  DFFPOSX1 DFFPOSX1_100 (.Q(regs_30__3_), .gnd(gnd), .vdd(vdd), .D(_761_), .CLK(clock_bf2__1), );
  DFFPOSX1 DFFPOSX1_101 (.Q(regs_30__4_), .gnd(gnd), .vdd(vdd), .D(_762_), .CLK(clock_bf2__12), );
  DFFPOSX1 DFFPOSX1_102 (.Q(regs_30__5_), .gnd(gnd), .vdd(vdd), .D(_763_), .CLK(random_clk_bf3__401), );
  DFFPOSX1 DFFPOSX1_103 (.Q(regs_30__6_), .gnd(gnd), .vdd(vdd), .D(_764_), .CLK(random_clk_bf3__621), );
  DFFPOSX1 DFFPOSX1_104 (.Q(regs_30__7_), .gnd(gnd), .vdd(vdd), .D(_765_), .CLK(random_clk_bf3__841), );
  DFFPOSX1 DFFPOSX1_105 (.Q(regs_30__8_), .gnd(gnd), .vdd(vdd), .D(_766_), .CLK(random_clk_bf3__1061), );
  DFFPOSX1 DFFPOSX1_106 (.Q(regs_30__9_), .gnd(gnd), .vdd(vdd), .D(_767_), .CLK(random_clk_bf3__1281), );
  DFFPOSX1 DFFPOSX1_107 (.Q(regs_30__10_), .gnd(gnd), .vdd(vdd), .D(_737_), .CLK(random_clk_bf3__1501), );
  DFFPOSX1 DFFPOSX1_108 (.Q(regs_30__11_), .gnd(gnd), .vdd(vdd), .D(_738_), .CLK(random_clk_bf3__1721), );
  DFFPOSX1 DFFPOSX1_109 (.Q(regs_30__12_), .gnd(gnd), .vdd(vdd), .D(_739_), .CLK(random_clk_bf3__1), );
  DFFPOSX1 DFFPOSX1_110 (.Q(regs_30__13_), .gnd(gnd), .vdd(vdd), .D(_740_), .CLK(random_clk_bf3__201), );
  DFFPOSX1 DFFPOSX1_111 (.Q(regs_30__14_), .gnd(gnd), .vdd(vdd), .D(_741_), .CLK(random_clk_bf3__421), );
  DFFPOSX1 DFFPOSX1_112 (.Q(regs_30__15_), .gnd(gnd), .vdd(vdd), .D(_742_), .CLK(random_clk_bf3__641), );
  DFFPOSX1 DFFPOSX1_113 (.Q(regs_30__16_), .gnd(gnd), .vdd(vdd), .D(_743_), .CLK(random_clk_bf3__861), );
  DFFPOSX1 DFFPOSX1_114 (.Q(regs_30__17_), .gnd(gnd), .vdd(vdd), .D(_744_), .CLK(random_clk_bf3__1081), );
  DFFPOSX1 DFFPOSX1_115 (.Q(regs_30__18_), .gnd(gnd), .vdd(vdd), .D(_745_), .CLK(random_clk_bf3__1301), );
  DFFPOSX1 DFFPOSX1_116 (.Q(regs_30__19_), .gnd(gnd), .vdd(vdd), .D(_746_), .CLK(random_clk_bf3__1521), );
  DFFPOSX1 DFFPOSX1_117 (.Q(regs_30__20_), .gnd(gnd), .vdd(vdd), .D(_748_), .CLK(random_clk_bf3__1741), );
  DFFPOSX1 DFFPOSX1_118 (.Q(regs_30__21_), .gnd(gnd), .vdd(vdd), .D(_749_), .CLK(random_clk_bf3__21), );
  DFFPOSX1 DFFPOSX1_119 (.Q(regs_30__22_), .gnd(gnd), .vdd(vdd), .D(_750_), .CLK(random_clk_bf3__221), );
  DFFPOSX1 DFFPOSX1_120 (.Q(regs_30__23_), .gnd(gnd), .vdd(vdd), .D(_751_), .CLK(random_clk_bf3__441), );
  DFFPOSX1 DFFPOSX1_121 (.Q(regs_30__24_), .gnd(gnd), .vdd(vdd), .D(_752_), .CLK(random_clk_bf3__661), );
  DFFPOSX1 DFFPOSX1_122 (.Q(regs_30__25_), .gnd(gnd), .vdd(vdd), .D(_753_), .CLK(random_clk_bf3__881), );
  DFFPOSX1 DFFPOSX1_123 (.Q(regs_30__26_), .gnd(gnd), .vdd(vdd), .D(_754_), .CLK(random_clk_bf3__1101), );
  DFFPOSX1 DFFPOSX1_124 (.Q(regs_30__27_), .gnd(gnd), .vdd(vdd), .D(_755_), .CLK(random_clk_bf3__1321), );
  DFFPOSX1 DFFPOSX1_125 (.Q(regs_30__28_), .gnd(gnd), .vdd(vdd), .D(_756_), .CLK(random_clk_bf3__1541), );
  DFFPOSX1 DFFPOSX1_126 (.Q(regs_30__29_), .gnd(gnd), .vdd(vdd), .D(_757_), .CLK(random_clk_bf3__1761), );
  DFFPOSX1 DFFPOSX1_127 (.Q(regs_30__30_), .gnd(gnd), .vdd(vdd), .D(_759_), .CLK(random_clk_bf3__41), );
  DFFPOSX1 DFFPOSX1_128 (.Q(regs_30__31_), .gnd(gnd), .vdd(vdd), .D(_760_), .CLK(random_clk_bf3__241), );
  DFFPOSX1 DFFPOSX1_129 (.Q(regs_29__0_), .gnd(gnd), .vdd(vdd), .D(_672_), .CLK(random_clk_bf3__461), );
  DFFPOSX1 DFFPOSX1_130 (.Q(regs_29__1_), .gnd(gnd), .vdd(vdd), .D(_683_), .CLK(random_clk_bf3__681), );
  DFFPOSX1 DFFPOSX1_131 (.Q(regs_29__2_), .gnd(gnd), .vdd(vdd), .D(_694_), .CLK(random_clk_bf3__901), );
  DFFPOSX1 DFFPOSX1_132 (.Q(regs_29__3_), .gnd(gnd), .vdd(vdd), .D(_697_), .CLK(random_clk_bf3__1121), );
  DFFPOSX1 DFFPOSX1_133 (.Q(regs_29__4_), .gnd(gnd), .vdd(vdd), .D(_698_), .CLK(random_clk_bf3__1341), );
  DFFPOSX1 DFFPOSX1_134 (.Q(regs_29__5_), .gnd(gnd), .vdd(vdd), .D(_699_), .CLK(random_clk_bf3__1561), );
  DFFPOSX1 DFFPOSX1_135 (.Q(regs_29__6_), .gnd(gnd), .vdd(vdd), .D(_700_), .CLK(random_clk_bf3__1781), );
  DFFPOSX1 DFFPOSX1_136 (.Q(regs_29__7_), .gnd(gnd), .vdd(vdd), .D(_701_), .CLK(random_clk_bf3__61), );
  DFFPOSX1 DFFPOSX1_137 (.Q(regs_29__8_), .gnd(gnd), .vdd(vdd), .D(_702_), .CLK(random_clk_bf3__261), );
  DFFPOSX1 DFFPOSX1_138 (.Q(regs_29__9_), .gnd(gnd), .vdd(vdd), .D(_703_), .CLK(random_clk_bf3__481), );
  DFFPOSX1 DFFPOSX1_139 (.Q(regs_29__10_), .gnd(gnd), .vdd(vdd), .D(_673_), .CLK(random_clk_bf3__701), );
  DFFPOSX1 DFFPOSX1_140 (.Q(regs_29__11_), .gnd(gnd), .vdd(vdd), .D(_674_), .CLK(random_clk_bf3__921), );
  DFFPOSX1 DFFPOSX1_141 (.Q(regs_29__12_), .gnd(gnd), .vdd(vdd), .D(_675_), .CLK(random_clk_bf3__1141), );
  DFFPOSX1 DFFPOSX1_142 (.Q(regs_29__13_), .gnd(gnd), .vdd(vdd), .D(_676_), .CLK(random_clk_bf3__1361), );
  DFFPOSX1 DFFPOSX1_143 (.Q(regs_29__14_), .gnd(gnd), .vdd(vdd), .D(_677_), .CLK(random_clk_bf3__1581), );
  DFFPOSX1 DFFPOSX1_144 (.Q(regs_29__15_), .gnd(gnd), .vdd(vdd), .D(_678_), .CLK(random_clk_bf3__1801), );
  DFFPOSX1 DFFPOSX1_145 (.Q(regs_29__16_), .gnd(gnd), .vdd(vdd), .D(_679_), .CLK(random_clk_bf3__81), );
  DFFPOSX1 DFFPOSX1_146 (.Q(regs_29__17_), .gnd(gnd), .vdd(vdd), .D(_680_), .CLK(random_clk_bf3__281), );
  DFFPOSX1 DFFPOSX1_147 (.Q(regs_29__18_), .gnd(gnd), .vdd(vdd), .D(_681_), .CLK(random_clk_bf3__501), );
  DFFPOSX1 DFFPOSX1_148 (.Q(regs_29__19_), .gnd(gnd), .vdd(vdd), .D(_682_), .CLK(random_clk_bf3__721), );
  DFFPOSX1 DFFPOSX1_149 (.Q(regs_29__20_), .gnd(gnd), .vdd(vdd), .D(_684_), .CLK(random_clk_bf3__941), );
  DFFPOSX1 DFFPOSX1_150 (.Q(regs_29__21_), .gnd(gnd), .vdd(vdd), .D(_685_), .CLK(random_clk_bf3__1161), );
  DFFPOSX1 DFFPOSX1_151 (.Q(regs_29__22_), .gnd(gnd), .vdd(vdd), .D(_686_), .CLK(random_clk_bf3__1381), );
  DFFPOSX1 DFFPOSX1_152 (.Q(regs_29__23_), .gnd(gnd), .vdd(vdd), .D(_687_), .CLK(random_clk_bf3__1601), );
  DFFPOSX1 DFFPOSX1_153 (.Q(regs_29__24_), .gnd(gnd), .vdd(vdd), .D(_688_), .CLK(random_clk_bf3__1821), );
  DFFPOSX1 DFFPOSX1_154 (.Q(regs_29__25_), .gnd(gnd), .vdd(vdd), .D(_689_), .CLK(random_clk_bf3__101), );
  DFFPOSX1 DFFPOSX1_155 (.Q(regs_29__26_), .gnd(gnd), .vdd(vdd), .D(_690_), .CLK(random_clk_bf3__301), );
  DFFPOSX1 DFFPOSX1_156 (.Q(regs_29__27_), .gnd(gnd), .vdd(vdd), .D(_691_), .CLK(random_clk_bf3__521), );
  DFFPOSX1 DFFPOSX1_157 (.Q(regs_29__28_), .gnd(gnd), .vdd(vdd), .D(_692_), .CLK(random_clk_bf3__741), );
  DFFPOSX1 DFFPOSX1_158 (.Q(regs_29__29_), .gnd(gnd), .vdd(vdd), .D(_693_), .CLK(random_clk_bf3__961), );
  DFFPOSX1 DFFPOSX1_159 (.Q(regs_29__30_), .gnd(gnd), .vdd(vdd), .D(_695_), .CLK(random_clk_bf3__1181), );
  DFFPOSX1 DFFPOSX1_160 (.Q(regs_29__31_), .gnd(gnd), .vdd(vdd), .D(_696_), .CLK(random_clk_bf3__1401), );
  DFFPOSX1 DFFPOSX1_161 (.Q(regs_27__0_), .gnd(gnd), .vdd(vdd), .D(_608_), .CLK(random_clk_bf3__1621), );
  DFFPOSX1 DFFPOSX1_162 (.Q(regs_27__1_), .gnd(gnd), .vdd(vdd), .D(_619_), .CLK(random_clk_bf3__1841), );
  DFFPOSX1 DFFPOSX1_163 (.Q(regs_27__2_), .gnd(gnd), .vdd(vdd), .D(_630_), .CLK(random_clk_bf3__121), );
  DFFPOSX1 DFFPOSX1_164 (.Q(regs_27__3_), .gnd(gnd), .vdd(vdd), .D(_633_), .CLK(random_clk_bf3__321), );
  DFFPOSX1 DFFPOSX1_165 (.Q(regs_27__4_), .gnd(gnd), .vdd(vdd), .D(_634_), .CLK(random_clk_bf3__541), );
  DFFPOSX1 DFFPOSX1_166 (.Q(regs_27__5_), .gnd(gnd), .vdd(vdd), .D(_635_), .CLK(random_clk_bf3__761), );
  DFFPOSX1 DFFPOSX1_167 (.Q(regs_27__6_), .gnd(gnd), .vdd(vdd), .D(_636_), .CLK(random_clk_bf3__981), );
  DFFPOSX1 DFFPOSX1_168 (.Q(regs_27__7_), .gnd(gnd), .vdd(vdd), .D(_637_), .CLK(random_clk_bf3__1201), );
  DFFPOSX1 DFFPOSX1_169 (.Q(regs_27__8_), .gnd(gnd), .vdd(vdd), .D(_638_), .CLK(random_clk_bf3__1421), );
  DFFPOSX1 DFFPOSX1_170 (.Q(regs_27__9_), .gnd(gnd), .vdd(vdd), .D(_639_), .CLK(random_clk_bf3__1641), );
  DFFPOSX1 DFFPOSX1_171 (.Q(regs_27__10_), .gnd(gnd), .vdd(vdd), .D(_609_), .CLK(random_clk_bf3__1861), );
  DFFPOSX1 DFFPOSX1_172 (.Q(regs_27__11_), .gnd(gnd), .vdd(vdd), .D(_610_), .CLK(random_clk_bf3__141), );
  DFFPOSX1 DFFPOSX1_173 (.Q(regs_27__12_), .gnd(gnd), .vdd(vdd), .D(_611_), .CLK(random_clk_bf3__341), );
  DFFPOSX1 DFFPOSX1_174 (.Q(regs_27__13_), .gnd(gnd), .vdd(vdd), .D(_612_), .CLK(random_clk_bf3__561), );
  DFFPOSX1 DFFPOSX1_175 (.Q(regs_27__14_), .gnd(gnd), .vdd(vdd), .D(_613_), .CLK(random_clk_bf3__781), );
  DFFPOSX1 DFFPOSX1_176 (.Q(regs_27__15_), .gnd(gnd), .vdd(vdd), .D(_614_), .CLK(random_clk_bf3__1001), );
  DFFPOSX1 DFFPOSX1_177 (.Q(regs_27__16_), .gnd(gnd), .vdd(vdd), .D(_615_), .CLK(random_clk_bf3__1221), );
  DFFPOSX1 DFFPOSX1_178 (.Q(regs_27__17_), .gnd(gnd), .vdd(vdd), .D(_616_), .CLK(random_clk_bf3__1441), );
  DFFPOSX1 DFFPOSX1_179 (.Q(regs_27__18_), .gnd(gnd), .vdd(vdd), .D(_617_), .CLK(random_clk_bf3__1661), );
  DFFPOSX1 DFFPOSX1_180 (.Q(regs_27__19_), .gnd(gnd), .vdd(vdd), .D(_618_), .CLK(random_clk_bf3__1881), );
  DFFPOSX1 DFFPOSX1_181 (.Q(regs_27__20_), .gnd(gnd), .vdd(vdd), .D(_620_), .CLK(random_clk_bf3__161), );
  DFFPOSX1 DFFPOSX1_182 (.Q(regs_27__21_), .gnd(gnd), .vdd(vdd), .D(_621_), .CLK(random_clk_bf3__361), );
  DFFPOSX1 DFFPOSX1_183 (.Q(regs_27__22_), .gnd(gnd), .vdd(vdd), .D(_622_), .CLK(random_clk_bf3__581), );
  DFFPOSX1 DFFPOSX1_184 (.Q(regs_27__23_), .gnd(gnd), .vdd(vdd), .D(_623_), .CLK(random_clk_bf3__801), );
  DFFPOSX1 DFFPOSX1_185 (.Q(regs_27__24_), .gnd(gnd), .vdd(vdd), .D(_624_), .CLK(random_clk_bf3__1021), );
  DFFPOSX1 DFFPOSX1_186 (.Q(regs_27__25_), .gnd(gnd), .vdd(vdd), .D(_625_), .CLK(random_clk_bf3__1241), );
  DFFPOSX1 DFFPOSX1_187 (.Q(regs_27__26_), .gnd(gnd), .vdd(vdd), .D(_626_), .CLK(random_clk_bf3__1461), );
  DFFPOSX1 DFFPOSX1_188 (.Q(regs_27__27_), .gnd(gnd), .vdd(vdd), .D(_627_), .CLK(random_clk_bf3__1681), );
  DFFPOSX1 DFFPOSX1_189 (.Q(regs_27__28_), .gnd(gnd), .vdd(vdd), .D(_628_), .CLK(random_clk_bf3__1901), );
  DFFPOSX1 DFFPOSX1_190 (.Q(regs_27__29_), .gnd(gnd), .vdd(vdd), .D(_629_), .CLK(random_clk_bf3__181), );
  DFFPOSX1 DFFPOSX1_191 (.Q(regs_27__30_), .gnd(gnd), .vdd(vdd), .D(_631_), .CLK(random_clk_bf3__381), );
  DFFPOSX1 DFFPOSX1_192 (.Q(regs_27__31_), .gnd(gnd), .vdd(vdd), .D(_632_), .CLK(random_clk_bf3__601), );
  DFFPOSX1 DFFPOSX1_193 (.Q(regs_26__0_), .gnd(gnd), .vdd(vdd), .D(_576_), .CLK(random_clk_bf3__821), );
  DFFPOSX1 DFFPOSX1_194 (.Q(regs_26__1_), .gnd(gnd), .vdd(vdd), .D(_587_), .CLK(random_clk_bf3__1041), );
  DFFPOSX1 DFFPOSX1_195 (.Q(regs_26__2_), .gnd(gnd), .vdd(vdd), .D(_598_), .CLK(random_clk_bf3__1261), );
  DFFPOSX1 DFFPOSX1_196 (.Q(regs_26__3_), .gnd(gnd), .vdd(vdd), .D(_601_), .CLK(random_clk_bf3__1481), );
  DFFPOSX1 DFFPOSX1_197 (.Q(regs_26__4_), .gnd(gnd), .vdd(vdd), .D(_602_), .CLK(random_clk_bf3__1701), );
  DFFPOSX1 DFFPOSX1_198 (.Q(regs_26__5_), .gnd(gnd), .vdd(vdd), .D(_603_), .CLK(clock_bf2__23), );
  DFFPOSX1 DFFPOSX1_199 (.Q(regs_26__6_), .gnd(gnd), .vdd(vdd), .D(_604_), .CLK(clock_bf2__2), );
  DFFPOSX1 DFFPOSX1_200 (.Q(regs_26__7_), .gnd(gnd), .vdd(vdd), .D(_605_), .CLK(clock_bf2__13), );
  DFFPOSX1 DFFPOSX1_201 (.Q(regs_26__8_), .gnd(gnd), .vdd(vdd), .D(_606_), .CLK(random_clk_bf3__401), );
  DFFPOSX1 DFFPOSX1_202 (.Q(regs_26__9_), .gnd(gnd), .vdd(vdd), .D(_607_), .CLK(random_clk_bf3__621), );
  DFFPOSX1 DFFPOSX1_203 (.Q(regs_26__10_), .gnd(gnd), .vdd(vdd), .D(_577_), .CLK(random_clk_bf3__841), );
  DFFPOSX1 DFFPOSX1_204 (.Q(regs_26__11_), .gnd(gnd), .vdd(vdd), .D(_578_), .CLK(random_clk_bf3__1061), );
  DFFPOSX1 DFFPOSX1_205 (.Q(regs_26__12_), .gnd(gnd), .vdd(vdd), .D(_579_), .CLK(random_clk_bf3__1281), );
  DFFPOSX1 DFFPOSX1_206 (.Q(regs_26__13_), .gnd(gnd), .vdd(vdd), .D(_580_), .CLK(random_clk_bf3__1501), );
  DFFPOSX1 DFFPOSX1_207 (.Q(regs_26__14_), .gnd(gnd), .vdd(vdd), .D(_581_), .CLK(random_clk_bf3__1721), );
  DFFPOSX1 DFFPOSX1_208 (.Q(regs_26__15_), .gnd(gnd), .vdd(vdd), .D(_582_), .CLK(random_clk_bf3__1), );
  DFFPOSX1 DFFPOSX1_209 (.Q(regs_26__16_), .gnd(gnd), .vdd(vdd), .D(_583_), .CLK(random_clk_bf3__201), );
  DFFPOSX1 DFFPOSX1_210 (.Q(regs_26__17_), .gnd(gnd), .vdd(vdd), .D(_584_), .CLK(random_clk_bf3__421), );
  DFFPOSX1 DFFPOSX1_211 (.Q(regs_26__18_), .gnd(gnd), .vdd(vdd), .D(_585_), .CLK(random_clk_bf3__641), );
  DFFPOSX1 DFFPOSX1_212 (.Q(regs_26__19_), .gnd(gnd), .vdd(vdd), .D(_586_), .CLK(random_clk_bf3__861), );
  DFFPOSX1 DFFPOSX1_213 (.Q(regs_26__20_), .gnd(gnd), .vdd(vdd), .D(_588_), .CLK(random_clk_bf3__1081), );
  DFFPOSX1 DFFPOSX1_214 (.Q(regs_26__21_), .gnd(gnd), .vdd(vdd), .D(_589_), .CLK(random_clk_bf3__1301), );
  DFFPOSX1 DFFPOSX1_215 (.Q(regs_26__22_), .gnd(gnd), .vdd(vdd), .D(_590_), .CLK(random_clk_bf3__1521), );
  DFFPOSX1 DFFPOSX1_216 (.Q(regs_26__23_), .gnd(gnd), .vdd(vdd), .D(_591_), .CLK(random_clk_bf3__1741), );
  DFFPOSX1 DFFPOSX1_217 (.Q(regs_26__24_), .gnd(gnd), .vdd(vdd), .D(_592_), .CLK(random_clk_bf3__21), );
  DFFPOSX1 DFFPOSX1_218 (.Q(regs_26__25_), .gnd(gnd), .vdd(vdd), .D(_593_), .CLK(random_clk_bf3__221), );
  DFFPOSX1 DFFPOSX1_219 (.Q(regs_26__26_), .gnd(gnd), .vdd(vdd), .D(_594_), .CLK(random_clk_bf3__441), );
  DFFPOSX1 DFFPOSX1_220 (.Q(regs_26__27_), .gnd(gnd), .vdd(vdd), .D(_595_), .CLK(random_clk_bf3__661), );
  DFFPOSX1 DFFPOSX1_221 (.Q(regs_26__28_), .gnd(gnd), .vdd(vdd), .D(_596_), .CLK(random_clk_bf3__881), );
  DFFPOSX1 DFFPOSX1_222 (.Q(regs_26__29_), .gnd(gnd), .vdd(vdd), .D(_597_), .CLK(random_clk_bf3__1101), );
  DFFPOSX1 DFFPOSX1_223 (.Q(regs_26__30_), .gnd(gnd), .vdd(vdd), .D(_599_), .CLK(random_clk_bf3__1321), );
  DFFPOSX1 DFFPOSX1_224 (.Q(regs_26__31_), .gnd(gnd), .vdd(vdd), .D(_600_), .CLK(random_clk_bf3__1541), );
  DFFPOSX1 DFFPOSX1_225 (.Q(regs_25__0_), .gnd(gnd), .vdd(vdd), .D(_544_), .CLK(random_clk_bf3__1761), );
  DFFPOSX1 DFFPOSX1_226 (.Q(regs_25__1_), .gnd(gnd), .vdd(vdd), .D(_555_), .CLK(random_clk_bf3__41), );
  DFFPOSX1 DFFPOSX1_227 (.Q(regs_25__2_), .gnd(gnd), .vdd(vdd), .D(_566_), .CLK(random_clk_bf3__241), );
  DFFPOSX1 DFFPOSX1_228 (.Q(regs_25__3_), .gnd(gnd), .vdd(vdd), .D(_569_), .CLK(random_clk_bf3__461), );
  DFFPOSX1 DFFPOSX1_229 (.Q(regs_25__4_), .gnd(gnd), .vdd(vdd), .D(_570_), .CLK(random_clk_bf3__681), );
  DFFPOSX1 DFFPOSX1_230 (.Q(regs_25__5_), .gnd(gnd), .vdd(vdd), .D(_571_), .CLK(random_clk_bf3__901), );
  DFFPOSX1 DFFPOSX1_231 (.Q(regs_25__6_), .gnd(gnd), .vdd(vdd), .D(_572_), .CLK(random_clk_bf3__1121), );
  DFFPOSX1 DFFPOSX1_232 (.Q(regs_25__7_), .gnd(gnd), .vdd(vdd), .D(_573_), .CLK(random_clk_bf3__1341), );
  DFFPOSX1 DFFPOSX1_233 (.Q(regs_25__8_), .gnd(gnd), .vdd(vdd), .D(_574_), .CLK(random_clk_bf3__1561), );
  DFFPOSX1 DFFPOSX1_234 (.Q(regs_25__9_), .gnd(gnd), .vdd(vdd), .D(_575_), .CLK(random_clk_bf3__1781), );
  DFFPOSX1 DFFPOSX1_235 (.Q(regs_25__10_), .gnd(gnd), .vdd(vdd), .D(_545_), .CLK(random_clk_bf3__61), );
  DFFPOSX1 DFFPOSX1_236 (.Q(regs_25__11_), .gnd(gnd), .vdd(vdd), .D(_546_), .CLK(random_clk_bf3__261), );
  DFFPOSX1 DFFPOSX1_237 (.Q(regs_25__12_), .gnd(gnd), .vdd(vdd), .D(_547_), .CLK(random_clk_bf3__481), );
  DFFPOSX1 DFFPOSX1_238 (.Q(regs_25__13_), .gnd(gnd), .vdd(vdd), .D(_548_), .CLK(random_clk_bf3__701), );
  DFFPOSX1 DFFPOSX1_239 (.Q(regs_25__14_), .gnd(gnd), .vdd(vdd), .D(_549_), .CLK(random_clk_bf3__921), );
  DFFPOSX1 DFFPOSX1_240 (.Q(regs_25__15_), .gnd(gnd), .vdd(vdd), .D(_550_), .CLK(random_clk_bf3__1141), );
  DFFPOSX1 DFFPOSX1_241 (.Q(regs_25__16_), .gnd(gnd), .vdd(vdd), .D(_551_), .CLK(random_clk_bf3__1361), );
  DFFPOSX1 DFFPOSX1_242 (.Q(regs_25__17_), .gnd(gnd), .vdd(vdd), .D(_552_), .CLK(random_clk_bf3__1581), );
  DFFPOSX1 DFFPOSX1_243 (.Q(regs_25__18_), .gnd(gnd), .vdd(vdd), .D(_553_), .CLK(random_clk_bf3__1801), );
  DFFPOSX1 DFFPOSX1_244 (.Q(regs_25__19_), .gnd(gnd), .vdd(vdd), .D(_554_), .CLK(random_clk_bf3__81), );
  DFFPOSX1 DFFPOSX1_245 (.Q(regs_25__20_), .gnd(gnd), .vdd(vdd), .D(_556_), .CLK(random_clk_bf3__281), );
  DFFPOSX1 DFFPOSX1_246 (.Q(regs_25__21_), .gnd(gnd), .vdd(vdd), .D(_557_), .CLK(random_clk_bf3__501), );
  DFFPOSX1 DFFPOSX1_247 (.Q(regs_25__22_), .gnd(gnd), .vdd(vdd), .D(_558_), .CLK(random_clk_bf3__721), );
  DFFPOSX1 DFFPOSX1_248 (.Q(regs_25__23_), .gnd(gnd), .vdd(vdd), .D(_559_), .CLK(random_clk_bf3__941), );
  DFFPOSX1 DFFPOSX1_249 (.Q(regs_25__24_), .gnd(gnd), .vdd(vdd), .D(_560_), .CLK(random_clk_bf3__1161), );
  DFFPOSX1 DFFPOSX1_250 (.Q(regs_25__25_), .gnd(gnd), .vdd(vdd), .D(_561_), .CLK(random_clk_bf3__1381), );
  DFFPOSX1 DFFPOSX1_251 (.Q(regs_25__26_), .gnd(gnd), .vdd(vdd), .D(_562_), .CLK(random_clk_bf3__1601), );
  DFFPOSX1 DFFPOSX1_252 (.Q(regs_25__27_), .gnd(gnd), .vdd(vdd), .D(_563_), .CLK(random_clk_bf3__1821), );
  DFFPOSX1 DFFPOSX1_253 (.Q(regs_25__28_), .gnd(gnd), .vdd(vdd), .D(_564_), .CLK(random_clk_bf3__101), );
  DFFPOSX1 DFFPOSX1_254 (.Q(regs_25__29_), .gnd(gnd), .vdd(vdd), .D(_565_), .CLK(random_clk_bf3__301), );
  DFFPOSX1 DFFPOSX1_255 (.Q(regs_25__30_), .gnd(gnd), .vdd(vdd), .D(_567_), .CLK(random_clk_bf3__521), );
  DFFPOSX1 DFFPOSX1_256 (.Q(regs_25__31_), .gnd(gnd), .vdd(vdd), .D(_568_), .CLK(random_clk_bf3__741), );
  DFFPOSX1 DFFPOSX1_257 (.Q(regs_24__0_), .gnd(gnd), .vdd(vdd), .D(_512_), .CLK(random_clk_bf3__961), );
  DFFPOSX1 DFFPOSX1_258 (.Q(regs_24__1_), .gnd(gnd), .vdd(vdd), .D(_523_), .CLK(random_clk_bf3__1181), );
  DFFPOSX1 DFFPOSX1_259 (.Q(regs_24__2_), .gnd(gnd), .vdd(vdd), .D(_534_), .CLK(random_clk_bf3__1401), );
  DFFPOSX1 DFFPOSX1_260 (.Q(regs_24__3_), .gnd(gnd), .vdd(vdd), .D(_537_), .CLK(random_clk_bf3__1621), );
  DFFPOSX1 DFFPOSX1_261 (.Q(regs_24__4_), .gnd(gnd), .vdd(vdd), .D(_538_), .CLK(random_clk_bf3__1841), );
  DFFPOSX1 DFFPOSX1_262 (.Q(regs_24__5_), .gnd(gnd), .vdd(vdd), .D(_539_), .CLK(random_clk_bf3__121), );
  DFFPOSX1 DFFPOSX1_263 (.Q(regs_24__6_), .gnd(gnd), .vdd(vdd), .D(_540_), .CLK(random_clk_bf3__321), );
  DFFPOSX1 DFFPOSX1_264 (.Q(regs_24__7_), .gnd(gnd), .vdd(vdd), .D(_541_), .CLK(random_clk_bf3__541), );
  DFFPOSX1 DFFPOSX1_265 (.Q(regs_24__8_), .gnd(gnd), .vdd(vdd), .D(_542_), .CLK(random_clk_bf3__761), );
  DFFPOSX1 DFFPOSX1_266 (.Q(regs_24__9_), .gnd(gnd), .vdd(vdd), .D(_543_), .CLK(random_clk_bf3__981), );
  DFFPOSX1 DFFPOSX1_267 (.Q(regs_24__10_), .gnd(gnd), .vdd(vdd), .D(_513_), .CLK(random_clk_bf3__1201), );
  DFFPOSX1 DFFPOSX1_268 (.Q(regs_24__11_), .gnd(gnd), .vdd(vdd), .D(_514_), .CLK(random_clk_bf3__1421), );
  DFFPOSX1 DFFPOSX1_269 (.Q(regs_24__12_), .gnd(gnd), .vdd(vdd), .D(_515_), .CLK(random_clk_bf3__1641), );
  DFFPOSX1 DFFPOSX1_270 (.Q(regs_24__13_), .gnd(gnd), .vdd(vdd), .D(_516_), .CLK(random_clk_bf3__1861), );
  DFFPOSX1 DFFPOSX1_271 (.Q(regs_24__14_), .gnd(gnd), .vdd(vdd), .D(_517_), .CLK(random_clk_bf3__141), );
  DFFPOSX1 DFFPOSX1_272 (.Q(regs_24__15_), .gnd(gnd), .vdd(vdd), .D(_518_), .CLK(random_clk_bf3__341), );
  DFFPOSX1 DFFPOSX1_273 (.Q(regs_24__16_), .gnd(gnd), .vdd(vdd), .D(_519_), .CLK(random_clk_bf3__561), );
  DFFPOSX1 DFFPOSX1_274 (.Q(regs_24__17_), .gnd(gnd), .vdd(vdd), .D(_520_), .CLK(random_clk_bf3__781), );
  DFFPOSX1 DFFPOSX1_275 (.Q(regs_24__18_), .gnd(gnd), .vdd(vdd), .D(_521_), .CLK(random_clk_bf3__1001), );
  DFFPOSX1 DFFPOSX1_276 (.Q(regs_24__19_), .gnd(gnd), .vdd(vdd), .D(_522_), .CLK(random_clk_bf3__1221), );
  DFFPOSX1 DFFPOSX1_277 (.Q(regs_24__20_), .gnd(gnd), .vdd(vdd), .D(_524_), .CLK(random_clk_bf3__1441), );
  DFFPOSX1 DFFPOSX1_278 (.Q(regs_24__21_), .gnd(gnd), .vdd(vdd), .D(_525_), .CLK(random_clk_bf3__1661), );
  DFFPOSX1 DFFPOSX1_279 (.Q(regs_24__22_), .gnd(gnd), .vdd(vdd), .D(_526_), .CLK(random_clk_bf3__1881), );
  DFFPOSX1 DFFPOSX1_280 (.Q(regs_24__23_), .gnd(gnd), .vdd(vdd), .D(_527_), .CLK(random_clk_bf3__161), );
  DFFPOSX1 DFFPOSX1_281 (.Q(regs_24__24_), .gnd(gnd), .vdd(vdd), .D(_528_), .CLK(random_clk_bf3__361), );
  DFFPOSX1 DFFPOSX1_282 (.Q(regs_24__25_), .gnd(gnd), .vdd(vdd), .D(_529_), .CLK(random_clk_bf3__581), );
  DFFPOSX1 DFFPOSX1_283 (.Q(regs_24__26_), .gnd(gnd), .vdd(vdd), .D(_530_), .CLK(random_clk_bf3__801), );
  DFFPOSX1 DFFPOSX1_284 (.Q(regs_24__27_), .gnd(gnd), .vdd(vdd), .D(_531_), .CLK(random_clk_bf3__1021), );
  DFFPOSX1 DFFPOSX1_285 (.Q(regs_24__28_), .gnd(gnd), .vdd(vdd), .D(_532_), .CLK(random_clk_bf3__1241), );
  DFFPOSX1 DFFPOSX1_286 (.Q(regs_24__29_), .gnd(gnd), .vdd(vdd), .D(_533_), .CLK(random_clk_bf3__1461), );
  DFFPOSX1 DFFPOSX1_287 (.Q(regs_24__30_), .gnd(gnd), .vdd(vdd), .D(_535_), .CLK(random_clk_bf3__1681), );
  DFFPOSX1 DFFPOSX1_288 (.Q(regs_24__31_), .gnd(gnd), .vdd(vdd), .D(_536_), .CLK(random_clk_bf3__1901), );
  DFFPOSX1 DFFPOSX1_289 (.Q(regs_23__0_), .gnd(gnd), .vdd(vdd), .D(_480_), .CLK(random_clk_bf3__181), );
  DFFPOSX1 DFFPOSX1_290 (.Q(regs_23__1_), .gnd(gnd), .vdd(vdd), .D(_491_), .CLK(random_clk_bf3__381), );
  DFFPOSX1 DFFPOSX1_291 (.Q(regs_23__2_), .gnd(gnd), .vdd(vdd), .D(_502_), .CLK(random_clk_bf3__601), );
  DFFPOSX1 DFFPOSX1_292 (.Q(regs_23__3_), .gnd(gnd), .vdd(vdd), .D(_505_), .CLK(random_clk_bf3__821), );
  DFFPOSX1 DFFPOSX1_293 (.Q(regs_23__4_), .gnd(gnd), .vdd(vdd), .D(_506_), .CLK(random_clk_bf3__1041), );
  DFFPOSX1 DFFPOSX1_294 (.Q(regs_23__5_), .gnd(gnd), .vdd(vdd), .D(_507_), .CLK(random_clk_bf3__1261), );
  DFFPOSX1 DFFPOSX1_295 (.Q(regs_23__6_), .gnd(gnd), .vdd(vdd), .D(_508_), .CLK(random_clk_bf3__1481), );
  DFFPOSX1 DFFPOSX1_296 (.Q(regs_23__7_), .gnd(gnd), .vdd(vdd), .D(_509_), .CLK(random_clk_bf3__1701), );
  DFFPOSX1 DFFPOSX1_297 (.Q(regs_23__8_), .gnd(gnd), .vdd(vdd), .D(_510_), .CLK(clock_bf2__24), );
  DFFPOSX1 DFFPOSX1_298 (.Q(regs_23__9_), .gnd(gnd), .vdd(vdd), .D(_511_), .CLK(clock_bf2__3), );
  DFFPOSX1 DFFPOSX1_299 (.Q(regs_23__10_), .gnd(gnd), .vdd(vdd), .D(_481_), .CLK(clock_bf2__14), );
  DFFPOSX1 DFFPOSX1_300 (.Q(regs_23__11_), .gnd(gnd), .vdd(vdd), .D(_482_), .CLK(random_clk_bf3__401), );
  DFFPOSX1 DFFPOSX1_301 (.Q(regs_23__12_), .gnd(gnd), .vdd(vdd), .D(_483_), .CLK(random_clk_bf3__621), );
  DFFPOSX1 DFFPOSX1_302 (.Q(regs_23__13_), .gnd(gnd), .vdd(vdd), .D(_484_), .CLK(random_clk_bf3__841), );
  DFFPOSX1 DFFPOSX1_303 (.Q(regs_23__14_), .gnd(gnd), .vdd(vdd), .D(_485_), .CLK(random_clk_bf3__1061), );
  DFFPOSX1 DFFPOSX1_304 (.Q(regs_23__15_), .gnd(gnd), .vdd(vdd), .D(_486_), .CLK(random_clk_bf3__1281), );
  DFFPOSX1 DFFPOSX1_305 (.Q(regs_23__16_), .gnd(gnd), .vdd(vdd), .D(_487_), .CLK(random_clk_bf3__1501), );
  DFFPOSX1 DFFPOSX1_306 (.Q(regs_23__17_), .gnd(gnd), .vdd(vdd), .D(_488_), .CLK(random_clk_bf3__1721), );
  DFFPOSX1 DFFPOSX1_307 (.Q(regs_23__18_), .gnd(gnd), .vdd(vdd), .D(_489_), .CLK(random_clk_bf3__1), );
  DFFPOSX1 DFFPOSX1_308 (.Q(regs_23__19_), .gnd(gnd), .vdd(vdd), .D(_490_), .CLK(random_clk_bf3__201), );
  DFFPOSX1 DFFPOSX1_309 (.Q(regs_23__20_), .gnd(gnd), .vdd(vdd), .D(_492_), .CLK(random_clk_bf3__421), );
  DFFPOSX1 DFFPOSX1_310 (.Q(regs_23__21_), .gnd(gnd), .vdd(vdd), .D(_493_), .CLK(random_clk_bf3__641), );
  DFFPOSX1 DFFPOSX1_311 (.Q(regs_23__22_), .gnd(gnd), .vdd(vdd), .D(_494_), .CLK(random_clk_bf3__861), );
  DFFPOSX1 DFFPOSX1_312 (.Q(regs_23__23_), .gnd(gnd), .vdd(vdd), .D(_495_), .CLK(random_clk_bf3__1081), );
  DFFPOSX1 DFFPOSX1_313 (.Q(regs_23__24_), .gnd(gnd), .vdd(vdd), .D(_496_), .CLK(random_clk_bf3__1301), );
  DFFPOSX1 DFFPOSX1_314 (.Q(regs_23__25_), .gnd(gnd), .vdd(vdd), .D(_497_), .CLK(random_clk_bf3__1521), );
  DFFPOSX1 DFFPOSX1_315 (.Q(regs_23__26_), .gnd(gnd), .vdd(vdd), .D(_498_), .CLK(random_clk_bf3__1741), );
  DFFPOSX1 DFFPOSX1_316 (.Q(regs_23__27_), .gnd(gnd), .vdd(vdd), .D(_499_), .CLK(random_clk_bf3__21), );
  DFFPOSX1 DFFPOSX1_317 (.Q(regs_23__28_), .gnd(gnd), .vdd(vdd), .D(_500_), .CLK(random_clk_bf3__221), );
  DFFPOSX1 DFFPOSX1_318 (.Q(regs_23__29_), .gnd(gnd), .vdd(vdd), .D(_501_), .CLK(random_clk_bf3__441), );
  DFFPOSX1 DFFPOSX1_319 (.Q(regs_23__30_), .gnd(gnd), .vdd(vdd), .D(_503_), .CLK(random_clk_bf3__661), );
  DFFPOSX1 DFFPOSX1_320 (.Q(regs_23__31_), .gnd(gnd), .vdd(vdd), .D(_504_), .CLK(random_clk_bf3__881), );
  DFFPOSX1 DFFPOSX1_321 (.Q(regs_22__0_), .gnd(gnd), .vdd(vdd), .D(_448_), .CLK(random_clk_bf3__1101), );
  DFFPOSX1 DFFPOSX1_322 (.Q(regs_22__1_), .gnd(gnd), .vdd(vdd), .D(_459_), .CLK(random_clk_bf3__1321), );
  DFFPOSX1 DFFPOSX1_323 (.Q(regs_22__2_), .gnd(gnd), .vdd(vdd), .D(_470_), .CLK(random_clk_bf3__1541), );
  DFFPOSX1 DFFPOSX1_324 (.Q(regs_22__3_), .gnd(gnd), .vdd(vdd), .D(_473_), .CLK(random_clk_bf3__1761), );
  DFFPOSX1 DFFPOSX1_325 (.Q(regs_22__4_), .gnd(gnd), .vdd(vdd), .D(_474_), .CLK(random_clk_bf3__41), );
  DFFPOSX1 DFFPOSX1_326 (.Q(regs_22__5_), .gnd(gnd), .vdd(vdd), .D(_475_), .CLK(random_clk_bf3__241), );
  DFFPOSX1 DFFPOSX1_327 (.Q(regs_22__6_), .gnd(gnd), .vdd(vdd), .D(_476_), .CLK(random_clk_bf3__461), );
  DFFPOSX1 DFFPOSX1_328 (.Q(regs_22__7_), .gnd(gnd), .vdd(vdd), .D(_477_), .CLK(random_clk_bf3__681), );
  DFFPOSX1 DFFPOSX1_329 (.Q(regs_22__8_), .gnd(gnd), .vdd(vdd), .D(_478_), .CLK(random_clk_bf3__901), );
  DFFPOSX1 DFFPOSX1_330 (.Q(regs_22__9_), .gnd(gnd), .vdd(vdd), .D(_479_), .CLK(random_clk_bf3__1121), );
  DFFPOSX1 DFFPOSX1_331 (.Q(regs_22__10_), .gnd(gnd), .vdd(vdd), .D(_449_), .CLK(random_clk_bf3__1341), );
  DFFPOSX1 DFFPOSX1_332 (.Q(regs_22__11_), .gnd(gnd), .vdd(vdd), .D(_450_), .CLK(random_clk_bf3__1561), );
  DFFPOSX1 DFFPOSX1_333 (.Q(regs_22__12_), .gnd(gnd), .vdd(vdd), .D(_451_), .CLK(random_clk_bf3__1781), );
  DFFPOSX1 DFFPOSX1_334 (.Q(regs_22__13_), .gnd(gnd), .vdd(vdd), .D(_452_), .CLK(random_clk_bf3__61), );
  DFFPOSX1 DFFPOSX1_335 (.Q(regs_22__14_), .gnd(gnd), .vdd(vdd), .D(_453_), .CLK(random_clk_bf3__261), );
  DFFPOSX1 DFFPOSX1_336 (.Q(regs_22__15_), .gnd(gnd), .vdd(vdd), .D(_454_), .CLK(random_clk_bf3__481), );
  DFFPOSX1 DFFPOSX1_337 (.Q(regs_22__16_), .gnd(gnd), .vdd(vdd), .D(_455_), .CLK(random_clk_bf3__701), );
  DFFPOSX1 DFFPOSX1_338 (.Q(regs_22__17_), .gnd(gnd), .vdd(vdd), .D(_456_), .CLK(random_clk_bf3__921), );
  DFFPOSX1 DFFPOSX1_339 (.Q(regs_22__18_), .gnd(gnd), .vdd(vdd), .D(_457_), .CLK(random_clk_bf3__1141), );
  DFFPOSX1 DFFPOSX1_340 (.Q(regs_22__19_), .gnd(gnd), .vdd(vdd), .D(_458_), .CLK(random_clk_bf3__1361), );
  DFFPOSX1 DFFPOSX1_341 (.Q(regs_22__20_), .gnd(gnd), .vdd(vdd), .D(_460_), .CLK(random_clk_bf3__1581), );
  DFFPOSX1 DFFPOSX1_342 (.Q(regs_22__21_), .gnd(gnd), .vdd(vdd), .D(_461_), .CLK(random_clk_bf3__1801), );
  DFFPOSX1 DFFPOSX1_343 (.Q(regs_22__22_), .gnd(gnd), .vdd(vdd), .D(_462_), .CLK(random_clk_bf3__81), );
  DFFPOSX1 DFFPOSX1_344 (.gnd(gnd), .Q(regs_22__23_), .vdd(vdd), .CLK(random_clk_bf3__281), .D(_463_), );
  DFFPOSX1 DFFPOSX1_345 (.gnd(gnd), .Q(regs_22__24_), .vdd(vdd), .CLK(random_clk_bf3__501), .D(_464_), );
  DFFPOSX1 DFFPOSX1_346 (.gnd(gnd), .Q(regs_22__25_), .vdd(vdd), .CLK(random_clk_bf3__721), .D(_465_), );
  DFFPOSX1 DFFPOSX1_347 (.gnd(gnd), .Q(regs_22__26_), .vdd(vdd), .CLK(random_clk_bf3__941), .D(_466_), );
  DFFPOSX1 DFFPOSX1_348 (.gnd(gnd), .Q(regs_22__27_), .vdd(vdd), .CLK(random_clk_bf3__1161), .D(_467_), );
  DFFPOSX1 DFFPOSX1_349 (.gnd(gnd), .Q(regs_22__28_), .vdd(vdd), .CLK(random_clk_bf3__1381), .D(_468_), );
  DFFPOSX1 DFFPOSX1_350 (.gnd(gnd), .Q(regs_22__29_), .vdd(vdd), .CLK(random_clk_bf3__1601), .D(_469_), );
  DFFPOSX1 DFFPOSX1_351 (.gnd(gnd), .Q(regs_22__30_), .vdd(vdd), .CLK(random_clk_bf3__1821), .D(_471_), );
  DFFPOSX1 DFFPOSX1_352 (.gnd(gnd), .Q(regs_22__31_), .vdd(vdd), .CLK(random_clk_bf3__101), .D(_472_), );
  DFFPOSX1 DFFPOSX1_353 (.gnd(gnd), .Q(regs_20__0_), .vdd(vdd), .CLK(random_clk_bf3__301), .D(_384_), );
  DFFPOSX1 DFFPOSX1_354 (.gnd(gnd), .Q(regs_20__1_), .vdd(vdd), .CLK(random_clk_bf3__521), .D(_395_), );
  DFFPOSX1 DFFPOSX1_355 (.gnd(gnd), .Q(regs_20__2_), .vdd(vdd), .CLK(random_clk_bf3__741), .D(_406_), );
  DFFPOSX1 DFFPOSX1_356 (.gnd(gnd), .Q(regs_20__3_), .vdd(vdd), .CLK(random_clk_bf3__961), .D(_409_), );
  DFFPOSX1 DFFPOSX1_357 (.gnd(gnd), .Q(regs_20__4_), .vdd(vdd), .CLK(random_clk_bf3__1181), .D(_410_), );
  DFFPOSX1 DFFPOSX1_358 (.gnd(gnd), .Q(regs_20__5_), .vdd(vdd), .CLK(random_clk_bf3__1401), .D(_411_), );
  DFFPOSX1 DFFPOSX1_359 (.gnd(gnd), .Q(regs_20__6_), .vdd(vdd), .CLK(random_clk_bf3__1621), .D(_412_), );
  DFFPOSX1 DFFPOSX1_360 (.gnd(gnd), .Q(regs_20__7_), .vdd(vdd), .CLK(random_clk_bf3__1841), .D(_413_), );
  DFFPOSX1 DFFPOSX1_361 (.gnd(gnd), .Q(regs_20__8_), .vdd(vdd), .CLK(random_clk_bf3__121), .D(_414_), );
  DFFPOSX1 DFFPOSX1_362 (.gnd(gnd), .Q(regs_20__9_), .vdd(vdd), .CLK(random_clk_bf3__321), .D(_415_), );
  DFFPOSX1 DFFPOSX1_363 (.gnd(gnd), .Q(regs_20__10_), .vdd(vdd), .CLK(random_clk_bf3__541), .D(_385_), );
  DFFPOSX1 DFFPOSX1_364 (.gnd(gnd), .Q(regs_20__11_), .vdd(vdd), .CLK(random_clk_bf3__761), .D(_386_), );
  DFFPOSX1 DFFPOSX1_365 (.gnd(gnd), .Q(regs_20__12_), .vdd(vdd), .CLK(random_clk_bf3__981), .D(_387_), );
  DFFPOSX1 DFFPOSX1_366 (.gnd(gnd), .Q(regs_20__13_), .vdd(vdd), .CLK(random_clk_bf3__1201), .D(_388_), );
  DFFPOSX1 DFFPOSX1_367 (.gnd(gnd), .Q(regs_20__14_), .vdd(vdd), .CLK(random_clk_bf3__1421), .D(_389_), );
  DFFPOSX1 DFFPOSX1_368 (.gnd(gnd), .Q(regs_20__15_), .vdd(vdd), .CLK(random_clk_bf3__1641), .D(_390_), );
  DFFPOSX1 DFFPOSX1_369 (.gnd(gnd), .Q(regs_20__16_), .vdd(vdd), .CLK(random_clk_bf3__1861), .D(_391_), );
  DFFPOSX1 DFFPOSX1_370 (.gnd(gnd), .Q(regs_20__17_), .vdd(vdd), .CLK(random_clk_bf3__141), .D(_392_), );
  DFFPOSX1 DFFPOSX1_371 (.gnd(gnd), .Q(regs_20__18_), .vdd(vdd), .CLK(random_clk_bf3__341), .D(_393_), );
  DFFPOSX1 DFFPOSX1_372 (.gnd(gnd), .Q(regs_20__19_), .vdd(vdd), .CLK(random_clk_bf3__561), .D(_394_), );
  DFFPOSX1 DFFPOSX1_373 (.gnd(gnd), .Q(regs_20__20_), .vdd(vdd), .CLK(random_clk_bf3__781), .D(_396_), );
  DFFPOSX1 DFFPOSX1_374 (.gnd(gnd), .Q(regs_20__21_), .vdd(vdd), .CLK(random_clk_bf3__1001), .D(_397_), );
  DFFPOSX1 DFFPOSX1_375 (.gnd(gnd), .Q(regs_20__22_), .vdd(vdd), .CLK(random_clk_bf3__1221), .D(_398_), );
  DFFPOSX1 DFFPOSX1_376 (.gnd(gnd), .Q(regs_20__23_), .vdd(vdd), .CLK(random_clk_bf3__1441), .D(_399_), );
  DFFPOSX1 DFFPOSX1_377 (.gnd(gnd), .Q(regs_20__24_), .vdd(vdd), .CLK(random_clk_bf3__1661), .D(_400_), );
  DFFPOSX1 DFFPOSX1_378 (.gnd(gnd), .Q(regs_20__25_), .vdd(vdd), .CLK(random_clk_bf3__1881), .D(_401_), );
  DFFPOSX1 DFFPOSX1_379 (.gnd(gnd), .Q(regs_20__26_), .vdd(vdd), .CLK(random_clk_bf3__161), .D(_402_), );
  DFFPOSX1 DFFPOSX1_380 (.gnd(gnd), .Q(regs_20__27_), .vdd(vdd), .CLK(random_clk_bf3__361), .D(_403_), );
  DFFPOSX1 DFFPOSX1_381 (.gnd(gnd), .Q(regs_20__28_), .vdd(vdd), .CLK(random_clk_bf3__581), .D(_404_), );
  DFFPOSX1 DFFPOSX1_382 (.gnd(gnd), .Q(regs_20__29_), .vdd(vdd), .CLK(random_clk_bf3__801), .D(_405_), );
  DFFPOSX1 DFFPOSX1_383 (.gnd(gnd), .Q(regs_20__30_), .vdd(vdd), .CLK(random_clk_bf3__1021), .D(_407_), );
  DFFPOSX1 DFFPOSX1_384 (.gnd(gnd), .Q(regs_20__31_), .vdd(vdd), .CLK(random_clk_bf3__1241), .D(_408_), );
  DFFPOSX1 DFFPOSX1_385 (.gnd(gnd), .Q(regs_21__0_), .vdd(vdd), .CLK(random_clk_bf3__1461), .D(_416_), );
  DFFPOSX1 DFFPOSX1_386 (.gnd(gnd), .Q(regs_21__1_), .vdd(vdd), .CLK(random_clk_bf3__1681), .D(_427_), );
  DFFPOSX1 DFFPOSX1_387 (.gnd(gnd), .Q(regs_21__2_), .vdd(vdd), .CLK(random_clk_bf3__1901), .D(_438_), );
  DFFPOSX1 DFFPOSX1_388 (.gnd(gnd), .Q(regs_21__3_), .vdd(vdd), .CLK(random_clk_bf3__181), .D(_441_), );
  DFFPOSX1 DFFPOSX1_389 (.gnd(gnd), .Q(regs_21__4_), .vdd(vdd), .CLK(random_clk_bf3__381), .D(_442_), );
  DFFPOSX1 DFFPOSX1_390 (.gnd(gnd), .Q(regs_21__5_), .vdd(vdd), .CLK(random_clk_bf3__601), .D(_443_), );
  DFFPOSX1 DFFPOSX1_391 (.gnd(gnd), .Q(regs_21__6_), .vdd(vdd), .CLK(random_clk_bf3__821), .D(_444_), );
  DFFPOSX1 DFFPOSX1_392 (.gnd(gnd), .Q(regs_21__7_), .vdd(vdd), .CLK(random_clk_bf3__1041), .D(_445_), );
  DFFPOSX1 DFFPOSX1_393 (.gnd(gnd), .Q(regs_21__8_), .vdd(vdd), .CLK(random_clk_bf3__1261), .D(_446_), );
  DFFPOSX1 DFFPOSX1_394 (.gnd(gnd), .Q(regs_21__9_), .vdd(vdd), .CLK(random_clk_bf3__1481), .D(_447_), );
  DFFPOSX1 DFFPOSX1_395 (.gnd(gnd), .Q(regs_21__10_), .vdd(vdd), .CLK(random_clk_bf3__1701), .D(_417_), );
  DFFPOSX1 DFFPOSX1_396 (.gnd(gnd), .Q(regs_21__11_), .vdd(vdd), .CLK(clock_bf2__25), .D(_418_), );
  DFFPOSX1 DFFPOSX1_397 (.gnd(gnd), .Q(regs_21__12_), .vdd(vdd), .CLK(clock_bf2__4), .D(_419_), );
  DFFPOSX1 DFFPOSX1_398 (.gnd(gnd), .Q(regs_21__13_), .vdd(vdd), .CLK(clock_bf2__15), .D(_420_), );
  DFFPOSX1 DFFPOSX1_399 (.gnd(gnd), .Q(regs_21__14_), .vdd(vdd), .CLK(random_clk_bf3__401), .D(_421_), );
  DFFPOSX1 DFFPOSX1_400 (.gnd(gnd), .Q(regs_21__15_), .vdd(vdd), .CLK(random_clk_bf3__621), .D(_422_), );
  DFFPOSX1 DFFPOSX1_401 (.gnd(gnd), .Q(regs_21__16_), .vdd(vdd), .CLK(random_clk_bf3__841), .D(_423_), );
  DFFPOSX1 DFFPOSX1_402 (.gnd(gnd), .Q(regs_21__17_), .vdd(vdd), .CLK(random_clk_bf3__1061), .D(_424_), );
  DFFPOSX1 DFFPOSX1_403 (.gnd(gnd), .Q(regs_21__18_), .vdd(vdd), .CLK(random_clk_bf3__1281), .D(_425_), );
  DFFPOSX1 DFFPOSX1_404 (.gnd(gnd), .Q(regs_21__19_), .vdd(vdd), .CLK(random_clk_bf3__1501), .D(_426_), );
  DFFPOSX1 DFFPOSX1_405 (.gnd(gnd), .Q(regs_21__20_), .vdd(vdd), .CLK(random_clk_bf3__1721), .D(_428_), );
  DFFPOSX1 DFFPOSX1_406 (.gnd(gnd), .Q(regs_21__21_), .vdd(vdd), .CLK(random_clk_bf3__1), .D(_429_), );
  DFFPOSX1 DFFPOSX1_407 (.gnd(gnd), .Q(regs_21__22_), .vdd(vdd), .CLK(random_clk_bf3__201), .D(_430_), );
  DFFPOSX1 DFFPOSX1_408 (.gnd(gnd), .Q(regs_21__23_), .vdd(vdd), .CLK(random_clk_bf3__421), .D(_431_), );
  DFFPOSX1 DFFPOSX1_409 (.gnd(gnd), .Q(regs_21__24_), .vdd(vdd), .CLK(random_clk_bf3__641), .D(_432_), );
  DFFPOSX1 DFFPOSX1_410 (.gnd(gnd), .Q(regs_21__25_), .vdd(vdd), .CLK(random_clk_bf3__861), .D(_433_), );
  DFFPOSX1 DFFPOSX1_411 (.gnd(gnd), .Q(regs_21__26_), .vdd(vdd), .CLK(random_clk_bf3__1081), .D(_434_), );
  DFFPOSX1 DFFPOSX1_412 (.gnd(gnd), .Q(regs_21__27_), .vdd(vdd), .CLK(random_clk_bf3__1301), .D(_435_), );
  DFFPOSX1 DFFPOSX1_413 (.gnd(gnd), .Q(regs_21__28_), .vdd(vdd), .CLK(random_clk_bf3__1521), .D(_436_), );
  DFFPOSX1 DFFPOSX1_414 (.gnd(gnd), .Q(regs_21__29_), .vdd(vdd), .CLK(random_clk_bf3__1741), .D(_437_), );
  DFFPOSX1 DFFPOSX1_415 (.gnd(gnd), .Q(regs_21__30_), .vdd(vdd), .CLK(random_clk_bf3__21), .D(_439_), );
  DFFPOSX1 DFFPOSX1_416 (.gnd(gnd), .Q(regs_21__31_), .vdd(vdd), .CLK(random_clk_bf3__221), .D(_440_), );
  DFFPOSX1 DFFPOSX1_417 (.gnd(gnd), .Q(regs_19__0_), .vdd(vdd), .CLK(random_clk_bf3__441), .D(_320_), );
  DFFPOSX1 DFFPOSX1_418 (.gnd(gnd), .Q(regs_19__1_), .vdd(vdd), .CLK(random_clk_bf3__661), .D(_331_), );
  DFFPOSX1 DFFPOSX1_419 (.gnd(gnd), .Q(regs_19__2_), .vdd(vdd), .CLK(random_clk_bf3__881), .D(_342_), );
  DFFPOSX1 DFFPOSX1_420 (.gnd(gnd), .Q(regs_19__3_), .vdd(vdd), .CLK(random_clk_bf3__1101), .D(_345_), );
  DFFPOSX1 DFFPOSX1_421 (.gnd(gnd), .Q(regs_19__4_), .vdd(vdd), .CLK(random_clk_bf3__1321), .D(_346_), );
  DFFPOSX1 DFFPOSX1_422 (.gnd(gnd), .Q(regs_19__5_), .vdd(vdd), .CLK(random_clk_bf3__1541), .D(_347_), );
  DFFPOSX1 DFFPOSX1_423 (.gnd(gnd), .Q(regs_19__6_), .vdd(vdd), .CLK(random_clk_bf3__1761), .D(_348_), );
  DFFPOSX1 DFFPOSX1_424 (.gnd(gnd), .Q(regs_19__7_), .vdd(vdd), .CLK(random_clk_bf3__41), .D(_349_), );
  DFFPOSX1 DFFPOSX1_425 (.gnd(gnd), .Q(regs_19__8_), .vdd(vdd), .CLK(random_clk_bf3__241), .D(_350_), );
  DFFPOSX1 DFFPOSX1_426 (.gnd(gnd), .Q(regs_19__9_), .vdd(vdd), .CLK(random_clk_bf3__461), .D(_351_), );
  DFFPOSX1 DFFPOSX1_427 (.gnd(gnd), .Q(regs_19__10_), .vdd(vdd), .CLK(random_clk_bf3__681), .D(_321_), );
  DFFPOSX1 DFFPOSX1_428 (.gnd(gnd), .Q(regs_19__11_), .vdd(vdd), .CLK(random_clk_bf3__901), .D(_322_), );
  DFFPOSX1 DFFPOSX1_429 (.gnd(gnd), .Q(regs_19__12_), .vdd(vdd), .CLK(random_clk_bf3__1121), .D(_323_), );
  DFFPOSX1 DFFPOSX1_430 (.gnd(gnd), .Q(regs_19__13_), .vdd(vdd), .CLK(random_clk_bf3__1341), .D(_324_), );
  DFFPOSX1 DFFPOSX1_431 (.gnd(gnd), .Q(regs_19__14_), .vdd(vdd), .CLK(random_clk_bf3__1561), .D(_325_), );
  DFFPOSX1 DFFPOSX1_432 (.gnd(gnd), .Q(regs_19__15_), .vdd(vdd), .CLK(random_clk_bf3__1781), .D(_326_), );
  DFFPOSX1 DFFPOSX1_433 (.gnd(gnd), .Q(regs_19__16_), .vdd(vdd), .CLK(random_clk_bf3__61), .D(_327_), );
  DFFPOSX1 DFFPOSX1_434 (.gnd(gnd), .Q(regs_19__17_), .vdd(vdd), .CLK(random_clk_bf3__261), .D(_328_), );
  DFFPOSX1 DFFPOSX1_435 (.gnd(gnd), .Q(regs_19__18_), .vdd(vdd), .CLK(random_clk_bf3__481), .D(_329_), );
  DFFPOSX1 DFFPOSX1_436 (.gnd(gnd), .Q(regs_19__19_), .vdd(vdd), .CLK(random_clk_bf3__701), .D(_330_), );
  DFFPOSX1 DFFPOSX1_437 (.gnd(gnd), .Q(regs_19__20_), .vdd(vdd), .CLK(random_clk_bf3__921), .D(_332_), );
  DFFPOSX1 DFFPOSX1_438 (.gnd(gnd), .Q(regs_19__21_), .vdd(vdd), .CLK(random_clk_bf3__1141), .D(_333_), );
  DFFPOSX1 DFFPOSX1_439 (.gnd(gnd), .Q(regs_19__22_), .vdd(vdd), .CLK(random_clk_bf3__1361), .D(_334_), );
  DFFPOSX1 DFFPOSX1_440 (.gnd(gnd), .Q(regs_19__23_), .vdd(vdd), .CLK(random_clk_bf3__1581), .D(_335_), );
  DFFPOSX1 DFFPOSX1_441 (.gnd(gnd), .Q(regs_19__24_), .vdd(vdd), .CLK(random_clk_bf3__1801), .D(_336_), );
  DFFPOSX1 DFFPOSX1_442 (.gnd(gnd), .Q(regs_19__25_), .vdd(vdd), .CLK(random_clk_bf3__81), .D(_337_), );
  DFFPOSX1 DFFPOSX1_443 (.gnd(gnd), .Q(regs_19__26_), .vdd(vdd), .CLK(random_clk_bf3__281), .D(_338_), );
  DFFPOSX1 DFFPOSX1_444 (.gnd(gnd), .Q(regs_19__27_), .vdd(vdd), .CLK(random_clk_bf3__501), .D(_339_), );
  DFFPOSX1 DFFPOSX1_445 (.gnd(gnd), .Q(regs_19__28_), .vdd(vdd), .CLK(random_clk_bf3__721), .D(_340_), );
  DFFPOSX1 DFFPOSX1_446 (.gnd(gnd), .Q(regs_19__29_), .vdd(vdd), .CLK(random_clk_bf3__941), .D(_341_), );
  DFFPOSX1 DFFPOSX1_447 (.gnd(gnd), .Q(regs_19__30_), .vdd(vdd), .CLK(random_clk_bf3__1161), .D(_343_), );
  DFFPOSX1 DFFPOSX1_448 (.gnd(gnd), .Q(regs_19__31_), .vdd(vdd), .CLK(random_clk_bf3__1381), .D(_344_), );
  DFFPOSX1 DFFPOSX1_449 (.gnd(gnd), .Q(regs_18__0_), .vdd(vdd), .CLK(random_clk_bf3__1601), .D(_288_), );
  DFFPOSX1 DFFPOSX1_450 (.gnd(gnd), .Q(regs_18__1_), .vdd(vdd), .CLK(random_clk_bf3__1821), .D(_299_), );
  DFFPOSX1 DFFPOSX1_451 (.gnd(gnd), .Q(regs_18__2_), .vdd(vdd), .CLK(random_clk_bf3__101), .D(_310_), );
  DFFPOSX1 DFFPOSX1_452 (.gnd(gnd), .Q(regs_18__3_), .vdd(vdd), .CLK(random_clk_bf3__301), .D(_313_), );
  DFFPOSX1 DFFPOSX1_453 (.gnd(gnd), .Q(regs_18__4_), .vdd(vdd), .CLK(random_clk_bf3__521), .D(_314_), );
  DFFPOSX1 DFFPOSX1_454 (.gnd(gnd), .Q(regs_18__5_), .vdd(vdd), .CLK(random_clk_bf3__741), .D(_315_), );
  DFFPOSX1 DFFPOSX1_455 (.gnd(gnd), .Q(regs_18__6_), .vdd(vdd), .CLK(random_clk_bf3__961), .D(_316_), );
  DFFPOSX1 DFFPOSX1_456 (.gnd(gnd), .Q(regs_18__7_), .vdd(vdd), .CLK(random_clk_bf3__1181), .D(_317_), );
  DFFPOSX1 DFFPOSX1_457 (.gnd(gnd), .Q(regs_18__8_), .vdd(vdd), .CLK(random_clk_bf3__1401), .D(_318_), );
  DFFPOSX1 DFFPOSX1_458 (.gnd(gnd), .Q(regs_18__9_), .vdd(vdd), .CLK(random_clk_bf3__1621), .D(_319_), );
  DFFPOSX1 DFFPOSX1_459 (.gnd(gnd), .Q(regs_18__10_), .vdd(vdd), .CLK(random_clk_bf3__1841), .D(_289_), );
  DFFPOSX1 DFFPOSX1_460 (.gnd(gnd), .Q(regs_18__11_), .vdd(vdd), .CLK(random_clk_bf3__121), .D(_290_), );
  DFFPOSX1 DFFPOSX1_461 (.gnd(gnd), .Q(regs_18__12_), .vdd(vdd), .CLK(random_clk_bf3__321), .D(_291_), );
  DFFPOSX1 DFFPOSX1_462 (.gnd(gnd), .Q(regs_18__13_), .vdd(vdd), .CLK(random_clk_bf3__541), .D(_292_), );
  DFFPOSX1 DFFPOSX1_463 (.gnd(gnd), .Q(regs_18__14_), .vdd(vdd), .CLK(random_clk_bf3__761), .D(_293_), );
  DFFPOSX1 DFFPOSX1_464 (.gnd(gnd), .Q(regs_18__15_), .vdd(vdd), .CLK(random_clk_bf3__981), .D(_294_), );
  DFFPOSX1 DFFPOSX1_465 (.gnd(gnd), .Q(regs_18__16_), .vdd(vdd), .CLK(random_clk_bf3__1201), .D(_295_), );
  DFFPOSX1 DFFPOSX1_466 (.gnd(gnd), .Q(regs_18__17_), .vdd(vdd), .CLK(random_clk_bf3__1421), .D(_296_), );
  DFFPOSX1 DFFPOSX1_467 (.gnd(gnd), .Q(regs_18__18_), .vdd(vdd), .CLK(random_clk_bf3__1641), .D(_297_), );
  DFFPOSX1 DFFPOSX1_468 (.gnd(gnd), .Q(regs_18__19_), .vdd(vdd), .CLK(random_clk_bf3__1861), .D(_298_), );
  DFFPOSX1 DFFPOSX1_469 (.gnd(gnd), .Q(regs_18__20_), .vdd(vdd), .CLK(random_clk_bf3__141), .D(_300_), );
  DFFPOSX1 DFFPOSX1_470 (.gnd(gnd), .Q(regs_18__21_), .vdd(vdd), .CLK(random_clk_bf3__341), .D(_301_), );
  DFFPOSX1 DFFPOSX1_471 (.gnd(gnd), .Q(regs_18__22_), .vdd(vdd), .CLK(random_clk_bf3__561), .D(_302_), );
  DFFPOSX1 DFFPOSX1_472 (.gnd(gnd), .Q(regs_18__23_), .vdd(vdd), .CLK(random_clk_bf3__781), .D(_303_), );
  DFFPOSX1 DFFPOSX1_473 (.gnd(gnd), .Q(regs_18__24_), .vdd(vdd), .CLK(random_clk_bf3__1001), .D(_304_), );
  DFFPOSX1 DFFPOSX1_474 (.gnd(gnd), .Q(regs_18__25_), .vdd(vdd), .CLK(random_clk_bf3__1221), .D(_305_), );
  DFFPOSX1 DFFPOSX1_475 (.gnd(gnd), .Q(regs_18__26_), .vdd(vdd), .CLK(random_clk_bf3__1441), .D(_306_), );
  DFFPOSX1 DFFPOSX1_476 (.gnd(gnd), .Q(regs_18__27_), .vdd(vdd), .CLK(random_clk_bf3__1661), .D(_307_), );
  DFFPOSX1 DFFPOSX1_477 (.gnd(gnd), .Q(regs_18__28_), .vdd(vdd), .CLK(random_clk_bf3__1881), .D(_308_), );
  DFFPOSX1 DFFPOSX1_478 (.gnd(gnd), .Q(regs_18__29_), .vdd(vdd), .CLK(random_clk_bf3__161), .D(_309_), );
  DFFPOSX1 DFFPOSX1_479 (.gnd(gnd), .Q(regs_18__30_), .vdd(vdd), .CLK(random_clk_bf3__361), .D(_311_), );
  DFFPOSX1 DFFPOSX1_480 (.gnd(gnd), .Q(regs_18__31_), .vdd(vdd), .CLK(random_clk_bf3__581), .D(_312_), );
  DFFPOSX1 DFFPOSX1_481 (.gnd(gnd), .Q(regs_17__0_), .vdd(vdd), .CLK(random_clk_bf3__801), .D(_256_), );
  DFFPOSX1 DFFPOSX1_482 (.gnd(gnd), .Q(regs_17__1_), .vdd(vdd), .CLK(random_clk_bf3__1021), .D(_267_), );
  DFFPOSX1 DFFPOSX1_483 (.gnd(gnd), .Q(regs_17__2_), .vdd(vdd), .CLK(random_clk_bf3__1241), .D(_278_), );
  DFFPOSX1 DFFPOSX1_484 (.gnd(gnd), .Q(regs_17__3_), .vdd(vdd), .CLK(random_clk_bf3__1461), .D(_281_), );
  DFFPOSX1 DFFPOSX1_485 (.gnd(gnd), .Q(regs_17__4_), .vdd(vdd), .CLK(random_clk_bf3__1681), .D(_282_), );
  DFFPOSX1 DFFPOSX1_486 (.gnd(gnd), .Q(regs_17__5_), .vdd(vdd), .CLK(random_clk_bf3__1901), .D(_283_), );
  DFFPOSX1 DFFPOSX1_487 (.gnd(gnd), .Q(regs_17__6_), .vdd(vdd), .CLK(random_clk_bf3__181), .D(_284_), );
  DFFPOSX1 DFFPOSX1_488 (.gnd(gnd), .Q(regs_17__7_), .vdd(vdd), .CLK(random_clk_bf3__381), .D(_285_), );
  DFFPOSX1 DFFPOSX1_489 (.gnd(gnd), .Q(regs_17__8_), .vdd(vdd), .CLK(random_clk_bf3__601), .D(_286_), );
  DFFPOSX1 DFFPOSX1_490 (.gnd(gnd), .Q(regs_17__9_), .vdd(vdd), .CLK(random_clk_bf3__821), .D(_287_), );
  DFFPOSX1 DFFPOSX1_491 (.gnd(gnd), .Q(regs_17__10_), .vdd(vdd), .CLK(random_clk_bf3__1041), .D(_257_), );
  DFFPOSX1 DFFPOSX1_492 (.gnd(gnd), .Q(regs_17__11_), .vdd(vdd), .CLK(random_clk_bf3__1261), .D(_258_), );
  DFFPOSX1 DFFPOSX1_493 (.gnd(gnd), .Q(regs_17__12_), .vdd(vdd), .CLK(random_clk_bf3__1481), .D(_259_), );
  DFFPOSX1 DFFPOSX1_494 (.gnd(gnd), .Q(regs_17__13_), .vdd(vdd), .CLK(random_clk_bf3__1701), .D(_260_), );
  DFFPOSX1 DFFPOSX1_495 (.gnd(gnd), .Q(regs_17__14_), .vdd(vdd), .CLK(clock_bf2__26), .D(_261_), );
  DFFPOSX1 DFFPOSX1_496 (.gnd(gnd), .Q(regs_17__15_), .vdd(vdd), .CLK(clock_bf2__5), .D(_262_), );
  DFFPOSX1 DFFPOSX1_497 (.gnd(gnd), .Q(regs_17__16_), .vdd(vdd), .CLK(clock_bf2__16), .D(_263_), );
  DFFPOSX1 DFFPOSX1_498 (.gnd(gnd), .Q(regs_17__17_), .vdd(vdd), .CLK(random_clk_bf3__402), .D(_264_), );
  DFFPOSX1 DFFPOSX1_499 (.gnd(gnd), .Q(regs_17__18_), .vdd(vdd), .CLK(random_clk_bf3__622), .D(_265_), );
  DFFPOSX1 DFFPOSX1_500 (.gnd(gnd), .Q(regs_17__19_), .vdd(vdd), .CLK(random_clk_bf3__842), .D(_266_), );
  DFFPOSX1 DFFPOSX1_501 (.gnd(gnd), .Q(regs_17__20_), .vdd(vdd), .CLK(random_clk_bf3__1062), .D(_268_), );
  DFFPOSX1 DFFPOSX1_502 (.gnd(gnd), .Q(regs_17__21_), .vdd(vdd), .CLK(random_clk_bf3__1282), .D(_269_), );
  DFFPOSX1 DFFPOSX1_503 (.gnd(gnd), .Q(regs_17__22_), .vdd(vdd), .CLK(random_clk_bf3__1502), .D(_270_), );
  DFFPOSX1 DFFPOSX1_504 (.gnd(gnd), .Q(regs_17__23_), .vdd(vdd), .CLK(random_clk_bf3__1722), .D(_271_), );
  DFFPOSX1 DFFPOSX1_505 (.gnd(gnd), .Q(regs_17__24_), .vdd(vdd), .CLK(random_clk_bf3__2), .D(_272_), );
  DFFPOSX1 DFFPOSX1_506 (.gnd(gnd), .Q(regs_17__25_), .vdd(vdd), .CLK(random_clk_bf3__202), .D(_273_), );
  DFFPOSX1 DFFPOSX1_507 (.gnd(gnd), .Q(regs_17__26_), .vdd(vdd), .CLK(random_clk_bf3__422), .D(_274_), );
  DFFPOSX1 DFFPOSX1_508 (.gnd(gnd), .Q(regs_17__27_), .vdd(vdd), .CLK(random_clk_bf3__642), .D(_275_), );
  DFFPOSX1 DFFPOSX1_509 (.gnd(gnd), .Q(regs_17__28_), .vdd(vdd), .CLK(random_clk_bf3__862), .D(_276_), );
  DFFPOSX1 DFFPOSX1_510 (.gnd(gnd), .Q(regs_17__29_), .vdd(vdd), .CLK(random_clk_bf3__1082), .D(_277_), );
  DFFPOSX1 DFFPOSX1_511 (.gnd(gnd), .Q(regs_17__30_), .vdd(vdd), .CLK(random_clk_bf3__1302), .D(_279_), );
  DFFPOSX1 DFFPOSX1_512 (.gnd(gnd), .Q(regs_17__31_), .vdd(vdd), .CLK(random_clk_bf3__1522), .D(_280_), );
  DFFPOSX1 DFFPOSX1_513 (.gnd(gnd), .Q(regs_16__0_), .vdd(vdd), .CLK(random_clk_bf3__1742), .D(_224_), );
  DFFPOSX1 DFFPOSX1_514 (.gnd(gnd), .Q(regs_16__1_), .vdd(vdd), .CLK(random_clk_bf3__22), .D(_235_), );
  DFFPOSX1 DFFPOSX1_515 (.gnd(gnd), .Q(regs_16__2_), .vdd(vdd), .CLK(random_clk_bf3__222), .D(_246_), );
  DFFPOSX1 DFFPOSX1_516 (.gnd(gnd), .Q(regs_16__3_), .vdd(vdd), .CLK(random_clk_bf3__442), .D(_249_), );
  DFFPOSX1 DFFPOSX1_517 (.gnd(gnd), .Q(regs_16__4_), .vdd(vdd), .CLK(random_clk_bf3__662), .D(_250_), );
  DFFPOSX1 DFFPOSX1_518 (.gnd(gnd), .Q(regs_16__5_), .vdd(vdd), .CLK(random_clk_bf3__882), .D(_251_), );
  DFFPOSX1 DFFPOSX1_519 (.gnd(gnd), .Q(regs_16__6_), .vdd(vdd), .CLK(random_clk_bf3__1102), .D(_252_), );
  DFFPOSX1 DFFPOSX1_520 (.gnd(gnd), .Q(regs_16__7_), .vdd(vdd), .CLK(random_clk_bf3__1322), .D(_253_), );
  DFFPOSX1 DFFPOSX1_521 (.gnd(gnd), .Q(regs_16__8_), .vdd(vdd), .CLK(random_clk_bf3__1542), .D(_254_), );
  DFFPOSX1 DFFPOSX1_522 (.gnd(gnd), .Q(regs_16__9_), .vdd(vdd), .CLK(random_clk_bf3__1762), .D(_255_), );
  DFFPOSX1 DFFPOSX1_523 (.gnd(gnd), .Q(regs_16__10_), .vdd(vdd), .CLK(random_clk_bf3__42), .D(_225_), );
  DFFPOSX1 DFFPOSX1_524 (.gnd(gnd), .Q(regs_16__11_), .vdd(vdd), .CLK(random_clk_bf3__242), .D(_226_), );
  DFFPOSX1 DFFPOSX1_525 (.gnd(gnd), .Q(regs_16__12_), .vdd(vdd), .CLK(random_clk_bf3__462), .D(_227_), );
  DFFPOSX1 DFFPOSX1_526 (.gnd(gnd), .Q(regs_16__13_), .vdd(vdd), .CLK(random_clk_bf3__682), .D(_228_), );
  DFFPOSX1 DFFPOSX1_527 (.gnd(gnd), .Q(regs_16__14_), .vdd(vdd), .CLK(random_clk_bf3__902), .D(_229_), );
  DFFPOSX1 DFFPOSX1_528 (.gnd(gnd), .Q(regs_16__15_), .vdd(vdd), .CLK(random_clk_bf3__1122), .D(_230_), );
  DFFPOSX1 DFFPOSX1_529 (.gnd(gnd), .Q(regs_16__16_), .vdd(vdd), .CLK(random_clk_bf3__1342), .D(_231_), );
  DFFPOSX1 DFFPOSX1_530 (.gnd(gnd), .Q(regs_16__17_), .vdd(vdd), .CLK(random_clk_bf3__1562), .D(_232_), );
  DFFPOSX1 DFFPOSX1_531 (.gnd(gnd), .Q(regs_16__18_), .vdd(vdd), .CLK(random_clk_bf3__1782), .D(_233_), );
  DFFPOSX1 DFFPOSX1_532 (.gnd(gnd), .Q(regs_16__19_), .vdd(vdd), .CLK(random_clk_bf3__62), .D(_234_), );
  DFFPOSX1 DFFPOSX1_533 (.gnd(gnd), .Q(regs_16__20_), .vdd(vdd), .CLK(random_clk_bf3__262), .D(_236_), );
  DFFPOSX1 DFFPOSX1_534 (.gnd(gnd), .Q(regs_16__21_), .vdd(vdd), .CLK(random_clk_bf3__482), .D(_237_), );
  DFFPOSX1 DFFPOSX1_535 (.gnd(gnd), .Q(regs_16__22_), .vdd(vdd), .CLK(random_clk_bf3__702), .D(_238_), );
  DFFPOSX1 DFFPOSX1_536 (.gnd(gnd), .Q(regs_16__23_), .vdd(vdd), .CLK(random_clk_bf3__922), .D(_239_), );
  DFFPOSX1 DFFPOSX1_537 (.gnd(gnd), .Q(regs_16__24_), .vdd(vdd), .CLK(random_clk_bf3__1142), .D(_240_), );
  DFFPOSX1 DFFPOSX1_538 (.gnd(gnd), .Q(regs_16__25_), .vdd(vdd), .CLK(random_clk_bf3__1362), .D(_241_), );
  DFFPOSX1 DFFPOSX1_539 (.gnd(gnd), .Q(regs_16__26_), .vdd(vdd), .CLK(random_clk_bf3__1582), .D(_242_), );
  DFFPOSX1 DFFPOSX1_540 (.gnd(gnd), .Q(regs_16__27_), .vdd(vdd), .CLK(random_clk_bf3__1802), .D(_243_), );
  DFFPOSX1 DFFPOSX1_541 (.gnd(gnd), .Q(regs_16__28_), .vdd(vdd), .CLK(random_clk_bf3__82), .D(_244_), );
  DFFPOSX1 DFFPOSX1_542 (.gnd(gnd), .Q(regs_16__29_), .vdd(vdd), .CLK(random_clk_bf3__282), .D(_245_), );
  DFFPOSX1 DFFPOSX1_543 (.gnd(gnd), .Q(regs_16__30_), .vdd(vdd), .CLK(random_clk_bf3__502), .D(_247_), );
  DFFPOSX1 DFFPOSX1_544 (.gnd(gnd), .Q(regs_16__31_), .vdd(vdd), .CLK(random_clk_bf3__722), .D(_248_), );
  DFFPOSX1 DFFPOSX1_545 (.gnd(gnd), .Q(regs_15__0_), .vdd(vdd), .CLK(random_clk_bf3__942), .D(_192_), );
  DFFPOSX1 DFFPOSX1_546 (.gnd(gnd), .Q(regs_15__1_), .vdd(vdd), .CLK(random_clk_bf3__1162), .D(_203_), );
  DFFPOSX1 DFFPOSX1_547 (.gnd(gnd), .Q(regs_15__2_), .vdd(vdd), .CLK(random_clk_bf3__1382), .D(_214_), );
  DFFPOSX1 DFFPOSX1_548 (.gnd(gnd), .Q(regs_15__3_), .vdd(vdd), .CLK(random_clk_bf3__1602), .D(_217_), );
  DFFPOSX1 DFFPOSX1_549 (.gnd(gnd), .Q(regs_15__4_), .vdd(vdd), .CLK(random_clk_bf3__1822), .D(_218_), );
  DFFPOSX1 DFFPOSX1_550 (.gnd(gnd), .Q(regs_15__5_), .vdd(vdd), .CLK(random_clk_bf3__102), .D(_219_), );
  DFFPOSX1 DFFPOSX1_551 (.gnd(gnd), .Q(regs_15__6_), .vdd(vdd), .CLK(random_clk_bf3__302), .D(_220_), );
  DFFPOSX1 DFFPOSX1_552 (.gnd(gnd), .Q(regs_15__7_), .vdd(vdd), .CLK(random_clk_bf3__522), .D(_221_), );
  DFFPOSX1 DFFPOSX1_553 (.gnd(gnd), .Q(regs_15__8_), .vdd(vdd), .CLK(random_clk_bf3__742), .D(_222_), );
  DFFPOSX1 DFFPOSX1_554 (.gnd(gnd), .Q(regs_15__9_), .vdd(vdd), .CLK(random_clk_bf3__962), .D(_223_), );
  DFFPOSX1 DFFPOSX1_555 (.gnd(gnd), .Q(regs_15__10_), .vdd(vdd), .CLK(random_clk_bf3__1182), .D(_193_), );
  DFFPOSX1 DFFPOSX1_556 (.gnd(gnd), .Q(regs_15__11_), .vdd(vdd), .CLK(random_clk_bf3__1402), .D(_194_), );
  DFFPOSX1 DFFPOSX1_557 (.gnd(gnd), .Q(regs_15__12_), .vdd(vdd), .CLK(random_clk_bf3__1622), .D(_195_), );
  DFFPOSX1 DFFPOSX1_558 (.gnd(gnd), .Q(regs_15__13_), .vdd(vdd), .CLK(random_clk_bf3__1842), .D(_196_), );
  DFFPOSX1 DFFPOSX1_559 (.gnd(gnd), .Q(regs_15__14_), .vdd(vdd), .CLK(random_clk_bf3__122), .D(_197_), );
  DFFPOSX1 DFFPOSX1_560 (.gnd(gnd), .Q(regs_15__15_), .vdd(vdd), .CLK(random_clk_bf3__322), .D(_198_), );
  DFFPOSX1 DFFPOSX1_561 (.gnd(gnd), .Q(regs_15__16_), .vdd(vdd), .CLK(random_clk_bf3__542), .D(_199_), );
  DFFPOSX1 DFFPOSX1_562 (.gnd(gnd), .Q(regs_15__17_), .vdd(vdd), .CLK(random_clk_bf3__762), .D(_200_), );
  DFFPOSX1 DFFPOSX1_563 (.gnd(gnd), .Q(regs_15__18_), .vdd(vdd), .CLK(random_clk_bf3__982), .D(_201_), );
  DFFPOSX1 DFFPOSX1_564 (.gnd(gnd), .Q(regs_15__19_), .vdd(vdd), .CLK(random_clk_bf3__1202), .D(_202_), );
  DFFPOSX1 DFFPOSX1_565 (.gnd(gnd), .Q(regs_15__20_), .vdd(vdd), .CLK(random_clk_bf3__1422), .D(_204_), );
  DFFPOSX1 DFFPOSX1_566 (.gnd(gnd), .Q(regs_15__21_), .vdd(vdd), .CLK(random_clk_bf3__1642), .D(_205_), );
  DFFPOSX1 DFFPOSX1_567 (.gnd(gnd), .Q(regs_15__22_), .vdd(vdd), .CLK(random_clk_bf3__1862), .D(_206_), );
  DFFPOSX1 DFFPOSX1_568 (.gnd(gnd), .Q(regs_15__23_), .vdd(vdd), .CLK(random_clk_bf3__142), .D(_207_), );
  DFFPOSX1 DFFPOSX1_569 (.gnd(gnd), .Q(regs_15__24_), .vdd(vdd), .CLK(random_clk_bf3__342), .D(_208_), );
  DFFPOSX1 DFFPOSX1_570 (.gnd(gnd), .Q(regs_15__25_), .vdd(vdd), .CLK(random_clk_bf3__562), .D(_209_), );
  DFFPOSX1 DFFPOSX1_571 (.gnd(gnd), .Q(regs_15__26_), .vdd(vdd), .CLK(random_clk_bf3__782), .D(_210_), );
  DFFPOSX1 DFFPOSX1_572 (.gnd(gnd), .Q(regs_15__27_), .vdd(vdd), .CLK(random_clk_bf3__1002), .D(_211_), );
  DFFPOSX1 DFFPOSX1_573 (.gnd(gnd), .Q(regs_15__28_), .vdd(vdd), .CLK(random_clk_bf3__1222), .D(_212_), );
  DFFPOSX1 DFFPOSX1_574 (.gnd(gnd), .Q(regs_15__29_), .vdd(vdd), .CLK(random_clk_bf3__1442), .D(_213_), );
  DFFPOSX1 DFFPOSX1_575 (.gnd(gnd), .Q(regs_15__30_), .vdd(vdd), .CLK(random_clk_bf3__1662), .D(_215_), );
  DFFPOSX1 DFFPOSX1_576 (.gnd(gnd), .Q(regs_15__31_), .vdd(vdd), .CLK(random_clk_bf3__1882), .D(_216_), );
  DFFPOSX1 DFFPOSX1_577 (.gnd(gnd), .Q(regs_14__0_), .vdd(vdd), .CLK(random_clk_bf3__162), .D(_160_), );
  DFFPOSX1 DFFPOSX1_578 (.gnd(gnd), .Q(regs_14__1_), .vdd(vdd), .CLK(random_clk_bf3__362), .D(_171_), );
  DFFPOSX1 DFFPOSX1_579 (.gnd(gnd), .Q(regs_14__2_), .vdd(vdd), .CLK(random_clk_bf3__582), .D(_182_), );
  DFFPOSX1 DFFPOSX1_580 (.gnd(gnd), .Q(regs_14__3_), .vdd(vdd), .CLK(random_clk_bf3__802), .D(_185_), );
  DFFPOSX1 DFFPOSX1_581 (.gnd(gnd), .Q(regs_14__4_), .vdd(vdd), .CLK(random_clk_bf3__1022), .D(_186_), );
  DFFPOSX1 DFFPOSX1_582 (.gnd(gnd), .Q(regs_14__5_), .vdd(vdd), .CLK(random_clk_bf3__1242), .D(_187_), );
  DFFPOSX1 DFFPOSX1_583 (.gnd(gnd), .Q(regs_14__6_), .vdd(vdd), .CLK(random_clk_bf3__1462), .D(_188_), );
  DFFPOSX1 DFFPOSX1_584 (.gnd(gnd), .Q(regs_14__7_), .vdd(vdd), .CLK(random_clk_bf3__1682), .D(_189_), );
  DFFPOSX1 DFFPOSX1_585 (.gnd(gnd), .Q(regs_14__8_), .vdd(vdd), .CLK(random_clk_bf3__1902), .D(_190_), );
  DFFPOSX1 DFFPOSX1_586 (.gnd(gnd), .Q(regs_14__9_), .vdd(vdd), .CLK(random_clk_bf3__182), .D(_191_), );
  DFFPOSX1 DFFPOSX1_587 (.gnd(gnd), .Q(regs_14__10_), .vdd(vdd), .CLK(random_clk_bf3__382), .D(_161_), );
  DFFPOSX1 DFFPOSX1_588 (.gnd(gnd), .Q(regs_14__11_), .vdd(vdd), .CLK(random_clk_bf3__602), .D(_162_), );
  DFFPOSX1 DFFPOSX1_589 (.gnd(gnd), .Q(regs_14__12_), .vdd(vdd), .CLK(random_clk_bf3__822), .D(_163_), );
  DFFPOSX1 DFFPOSX1_590 (.gnd(gnd), .Q(regs_14__13_), .vdd(vdd), .CLK(random_clk_bf3__1042), .D(_164_), );
  DFFPOSX1 DFFPOSX1_591 (.gnd(gnd), .Q(regs_14__14_), .vdd(vdd), .CLK(random_clk_bf3__1262), .D(_165_), );
  DFFPOSX1 DFFPOSX1_592 (.gnd(gnd), .Q(regs_14__15_), .vdd(vdd), .CLK(random_clk_bf3__1482), .D(_166_), );
  DFFPOSX1 DFFPOSX1_593 (.gnd(gnd), .Q(regs_14__16_), .vdd(vdd), .CLK(random_clk_bf3__1702), .D(_167_), );
  DFFPOSX1 DFFPOSX1_594 (.gnd(gnd), .Q(regs_14__17_), .vdd(vdd), .CLK(clock_bf2__27), .D(_168_), );
  DFFPOSX1 DFFPOSX1_595 (.gnd(gnd), .Q(regs_14__18_), .vdd(vdd), .CLK(clock_bf2__6), .D(_169_), );
  DFFPOSX1 DFFPOSX1_596 (.gnd(gnd), .Q(regs_14__19_), .vdd(vdd), .CLK(clock_bf2__17), .D(_170_), );
  DFFPOSX1 DFFPOSX1_597 (.gnd(gnd), .Q(regs_14__20_), .vdd(vdd), .CLK(random_clk_bf3__402), .D(_172_), );
  DFFPOSX1 DFFPOSX1_598 (.gnd(gnd), .Q(regs_14__21_), .vdd(vdd), .CLK(random_clk_bf3__622), .D(_173_), );
  DFFPOSX1 DFFPOSX1_599 (.gnd(gnd), .Q(regs_14__22_), .vdd(vdd), .CLK(random_clk_bf3__842), .D(_174_), );
  DFFPOSX1 DFFPOSX1_600 (.gnd(gnd), .Q(regs_14__23_), .vdd(vdd), .CLK(random_clk_bf3__1062), .D(_175_), );
  DFFPOSX1 DFFPOSX1_601 (.gnd(gnd), .Q(regs_14__24_), .vdd(vdd), .CLK(random_clk_bf3__1282), .D(_176_), );
  DFFPOSX1 DFFPOSX1_602 (.gnd(gnd), .Q(regs_14__25_), .vdd(vdd), .CLK(random_clk_bf3__1502), .D(_177_), );
  DFFPOSX1 DFFPOSX1_603 (.gnd(gnd), .Q(regs_14__26_), .vdd(vdd), .CLK(random_clk_bf3__1722), .D(_178_), );
  DFFPOSX1 DFFPOSX1_604 (.gnd(gnd), .Q(regs_14__27_), .vdd(vdd), .CLK(random_clk_bf3__2), .D(_179_), );
  DFFPOSX1 DFFPOSX1_605 (.gnd(gnd), .Q(regs_14__28_), .vdd(vdd), .CLK(random_clk_bf3__202), .D(_180_), );
  DFFPOSX1 DFFPOSX1_606 (.gnd(gnd), .Q(regs_14__29_), .vdd(vdd), .CLK(random_clk_bf3__422), .D(_181_), );
  DFFPOSX1 DFFPOSX1_607 (.gnd(gnd), .Q(regs_14__30_), .vdd(vdd), .CLK(random_clk_bf3__642), .D(_183_), );
  DFFPOSX1 DFFPOSX1_608 (.gnd(gnd), .Q(regs_14__31_), .vdd(vdd), .CLK(random_clk_bf3__862), .D(_184_), );
  DFFPOSX1 DFFPOSX1_609 (.gnd(gnd), .Q(regs_13__0_), .vdd(vdd), .CLK(random_clk_bf3__1082), .D(_128_), );
  DFFPOSX1 DFFPOSX1_610 (.gnd(gnd), .Q(regs_13__1_), .vdd(vdd), .CLK(random_clk_bf3__1302), .D(_139_), );
  DFFPOSX1 DFFPOSX1_611 (.gnd(gnd), .Q(regs_13__2_), .vdd(vdd), .CLK(random_clk_bf3__1522), .D(_150_), );
  DFFPOSX1 DFFPOSX1_612 (.gnd(gnd), .Q(regs_13__3_), .vdd(vdd), .CLK(random_clk_bf3__1742), .D(_153_), );
  DFFPOSX1 DFFPOSX1_613 (.gnd(gnd), .Q(regs_13__4_), .vdd(vdd), .CLK(random_clk_bf3__22), .D(_154_), );
  DFFPOSX1 DFFPOSX1_614 (.gnd(gnd), .Q(regs_13__5_), .vdd(vdd), .CLK(random_clk_bf3__222), .D(_155_), );
  DFFPOSX1 DFFPOSX1_615 (.gnd(gnd), .Q(regs_13__6_), .vdd(vdd), .CLK(random_clk_bf3__442), .D(_156_), );
  DFFPOSX1 DFFPOSX1_616 (.gnd(gnd), .Q(regs_13__7_), .vdd(vdd), .CLK(random_clk_bf3__662), .D(_157_), );
  DFFPOSX1 DFFPOSX1_617 (.gnd(gnd), .Q(regs_13__8_), .vdd(vdd), .CLK(random_clk_bf3__882), .D(_158_), );
  DFFPOSX1 DFFPOSX1_618 (.gnd(gnd), .Q(regs_13__9_), .vdd(vdd), .CLK(random_clk_bf3__1102), .D(_159_), );
  DFFPOSX1 DFFPOSX1_619 (.gnd(gnd), .Q(regs_13__10_), .vdd(vdd), .CLK(random_clk_bf3__1322), .D(_129_), );
  DFFPOSX1 DFFPOSX1_620 (.gnd(gnd), .Q(regs_13__11_), .vdd(vdd), .CLK(random_clk_bf3__1542), .D(_130_), );
  DFFPOSX1 DFFPOSX1_621 (.gnd(gnd), .Q(regs_13__12_), .vdd(vdd), .CLK(random_clk_bf3__1762), .D(_131_), );
  DFFPOSX1 DFFPOSX1_622 (.gnd(gnd), .Q(regs_13__13_), .vdd(vdd), .CLK(random_clk_bf3__42), .D(_132_), );
  DFFPOSX1 DFFPOSX1_623 (.gnd(gnd), .Q(regs_13__14_), .vdd(vdd), .CLK(random_clk_bf3__242), .D(_133_), );
  DFFPOSX1 DFFPOSX1_624 (.gnd(gnd), .Q(regs_13__15_), .vdd(vdd), .CLK(random_clk_bf3__462), .D(_134_), );
  DFFPOSX1 DFFPOSX1_625 (.gnd(gnd), .Q(regs_13__16_), .vdd(vdd), .CLK(random_clk_bf3__682), .D(_135_), );
  DFFPOSX1 DFFPOSX1_626 (.gnd(gnd), .Q(regs_13__17_), .vdd(vdd), .CLK(random_clk_bf3__902), .D(_136_), );
  DFFPOSX1 DFFPOSX1_627 (.gnd(gnd), .Q(regs_13__18_), .vdd(vdd), .CLK(random_clk_bf3__1122), .D(_137_), );
  DFFPOSX1 DFFPOSX1_628 (.gnd(gnd), .Q(regs_13__19_), .vdd(vdd), .CLK(random_clk_bf3__1342), .D(_138_), );
  DFFPOSX1 DFFPOSX1_629 (.gnd(gnd), .Q(regs_13__20_), .vdd(vdd), .CLK(random_clk_bf3__1562), .D(_140_), );
  DFFPOSX1 DFFPOSX1_630 (.gnd(gnd), .Q(regs_13__21_), .vdd(vdd), .CLK(random_clk_bf3__1782), .D(_141_), );
  DFFPOSX1 DFFPOSX1_631 (.gnd(gnd), .Q(regs_13__22_), .vdd(vdd), .CLK(random_clk_bf3__62), .D(_142_), );
  DFFPOSX1 DFFPOSX1_632 (.gnd(gnd), .Q(regs_13__23_), .vdd(vdd), .CLK(random_clk_bf3__262), .D(_143_), );
  DFFPOSX1 DFFPOSX1_633 (.gnd(gnd), .Q(regs_13__24_), .vdd(vdd), .CLK(random_clk_bf3__482), .D(_144_), );
  DFFPOSX1 DFFPOSX1_634 (.gnd(gnd), .Q(regs_13__25_), .vdd(vdd), .CLK(random_clk_bf3__702), .D(_145_), );
  DFFPOSX1 DFFPOSX1_635 (.gnd(gnd), .Q(regs_13__26_), .vdd(vdd), .CLK(random_clk_bf3__922), .D(_146_), );
  DFFPOSX1 DFFPOSX1_636 (.gnd(gnd), .Q(regs_13__27_), .vdd(vdd), .CLK(random_clk_bf3__1142), .D(_147_), );
  DFFPOSX1 DFFPOSX1_637 (.gnd(gnd), .Q(regs_13__28_), .vdd(vdd), .CLK(random_clk_bf3__1362), .D(_148_), );
  DFFPOSX1 DFFPOSX1_638 (.gnd(gnd), .Q(regs_13__29_), .vdd(vdd), .CLK(random_clk_bf3__1582), .D(_149_), );
  DFFPOSX1 DFFPOSX1_639 (.gnd(gnd), .Q(regs_13__30_), .vdd(vdd), .CLK(random_clk_bf3__1802), .D(_151_), );
  DFFPOSX1 DFFPOSX1_640 (.gnd(gnd), .Q(regs_13__31_), .vdd(vdd), .CLK(random_clk_bf3__82), .D(_152_), );
  DFFPOSX1 DFFPOSX1_641 (.gnd(gnd), .Q(regs_11__0_), .vdd(vdd), .CLK(random_clk_bf3__282), .D(_64_), );
  DFFPOSX1 DFFPOSX1_642 (.gnd(gnd), .Q(regs_11__1_), .vdd(vdd), .CLK(random_clk_bf3__502), .D(_75_), );
  DFFPOSX1 DFFPOSX1_643 (.gnd(gnd), .Q(regs_11__2_), .vdd(vdd), .CLK(random_clk_bf3__722), .D(_86_), );
  DFFPOSX1 DFFPOSX1_644 (.gnd(gnd), .Q(regs_11__3_), .vdd(vdd), .CLK(random_clk_bf3__942), .D(_89_), );
  DFFPOSX1 DFFPOSX1_645 (.gnd(gnd), .Q(regs_11__4_), .vdd(vdd), .CLK(random_clk_bf3__1162), .D(_90_), );
  DFFPOSX1 DFFPOSX1_646 (.gnd(gnd), .Q(regs_11__5_), .vdd(vdd), .CLK(random_clk_bf3__1382), .D(_91_), );
  DFFPOSX1 DFFPOSX1_647 (.gnd(gnd), .Q(regs_11__6_), .vdd(vdd), .CLK(random_clk_bf3__1602), .D(_92_), );
  DFFPOSX1 DFFPOSX1_648 (.gnd(gnd), .Q(regs_11__7_), .vdd(vdd), .CLK(random_clk_bf3__1822), .D(_93_), );
  DFFPOSX1 DFFPOSX1_649 (.gnd(gnd), .Q(regs_11__8_), .vdd(vdd), .CLK(random_clk_bf3__102), .D(_94_), );
  DFFPOSX1 DFFPOSX1_650 (.gnd(gnd), .Q(regs_11__9_), .vdd(vdd), .CLK(random_clk_bf3__302), .D(_95_), );
  DFFPOSX1 DFFPOSX1_651 (.gnd(gnd), .Q(regs_11__10_), .vdd(vdd), .CLK(random_clk_bf3__522), .D(_65_), );
  DFFPOSX1 DFFPOSX1_652 (.gnd(gnd), .Q(regs_11__11_), .vdd(vdd), .CLK(random_clk_bf3__742), .D(_66_), );
  DFFPOSX1 DFFPOSX1_653 (.gnd(gnd), .Q(regs_11__12_), .vdd(vdd), .CLK(random_clk_bf3__962), .D(_67_), );
  DFFPOSX1 DFFPOSX1_654 (.gnd(gnd), .Q(regs_11__13_), .vdd(vdd), .CLK(random_clk_bf3__1182), .D(_68_), );
  DFFPOSX1 DFFPOSX1_655 (.gnd(gnd), .Q(regs_11__14_), .vdd(vdd), .CLK(random_clk_bf3__1402), .D(_69_), );
  DFFPOSX1 DFFPOSX1_656 (.gnd(gnd), .Q(regs_11__15_), .vdd(vdd), .CLK(random_clk_bf3__1622), .D(_70_), );
  DFFPOSX1 DFFPOSX1_657 (.gnd(gnd), .Q(regs_11__16_), .vdd(vdd), .CLK(random_clk_bf3__1842), .D(_71_), );
  DFFPOSX1 DFFPOSX1_658 (.gnd(gnd), .Q(regs_11__17_), .vdd(vdd), .CLK(random_clk_bf3__122), .D(_72_), );
  DFFPOSX1 DFFPOSX1_659 (.gnd(gnd), .Q(regs_11__18_), .vdd(vdd), .CLK(random_clk_bf3__322), .D(_73_), );
  DFFPOSX1 DFFPOSX1_660 (.gnd(gnd), .Q(regs_11__19_), .vdd(vdd), .CLK(random_clk_bf3__542), .D(_74_), );
  DFFPOSX1 DFFPOSX1_661 (.gnd(gnd), .Q(regs_11__20_), .vdd(vdd), .CLK(random_clk_bf3__762), .D(_76_), );
  DFFPOSX1 DFFPOSX1_662 (.gnd(gnd), .Q(regs_11__21_), .vdd(vdd), .CLK(random_clk_bf3__982), .D(_77_), );
  DFFPOSX1 DFFPOSX1_663 (.gnd(gnd), .Q(regs_11__22_), .vdd(vdd), .CLK(random_clk_bf3__1202), .D(_78_), );
  DFFPOSX1 DFFPOSX1_664 (.gnd(gnd), .Q(regs_11__23_), .vdd(vdd), .CLK(random_clk_bf3__1422), .D(_79_), );
  DFFPOSX1 DFFPOSX1_665 (.gnd(gnd), .Q(regs_11__24_), .vdd(vdd), .CLK(random_clk_bf3__1642), .D(_80_), );
  DFFPOSX1 DFFPOSX1_666 (.gnd(gnd), .Q(regs_11__25_), .vdd(vdd), .CLK(random_clk_bf3__1862), .D(_81_), );
  DFFPOSX1 DFFPOSX1_667 (.gnd(gnd), .Q(regs_11__26_), .vdd(vdd), .CLK(random_clk_bf3__142), .D(_82_), );
  DFFPOSX1 DFFPOSX1_668 (.gnd(gnd), .Q(regs_11__27_), .vdd(vdd), .CLK(random_clk_bf3__342), .D(_83_), );
  DFFPOSX1 DFFPOSX1_669 (.gnd(gnd), .Q(regs_11__28_), .vdd(vdd), .CLK(random_clk_bf3__562), .D(_84_), );
  DFFPOSX1 DFFPOSX1_670 (.gnd(gnd), .Q(regs_11__29_), .vdd(vdd), .CLK(random_clk_bf3__782), .D(_85_), );
  DFFPOSX1 DFFPOSX1_671 (.gnd(gnd), .Q(regs_11__30_), .vdd(vdd), .CLK(random_clk_bf3__1002), .D(_87_), );
  DFFPOSX1 DFFPOSX1_672 (.gnd(gnd), .Q(regs_11__31_), .vdd(vdd), .CLK(random_clk_bf3__1222), .D(_88_), );
  DFFPOSX1 DFFPOSX1_673 (.gnd(gnd), .Q(regs_12__0_), .vdd(vdd), .CLK(random_clk_bf3__1442), .D(_96_), );
  DFFPOSX1 DFFPOSX1_674 (.gnd(gnd), .Q(regs_12__1_), .vdd(vdd), .CLK(random_clk_bf3__1662), .D(_107_), );
  DFFPOSX1 DFFPOSX1_675 (.gnd(gnd), .Q(regs_12__2_), .vdd(vdd), .CLK(random_clk_bf3__1882), .D(_118_), );
  DFFPOSX1 DFFPOSX1_676 (.gnd(gnd), .Q(regs_12__3_), .vdd(vdd), .CLK(random_clk_bf3__162), .D(_121_), );
  DFFPOSX1 DFFPOSX1_677 (.gnd(gnd), .Q(regs_12__4_), .vdd(vdd), .CLK(random_clk_bf3__362), .D(_122_), );
  DFFPOSX1 DFFPOSX1_678 (.gnd(gnd), .Q(regs_12__5_), .vdd(vdd), .CLK(random_clk_bf3__582), .D(_123_), );
  DFFPOSX1 DFFPOSX1_679 (.gnd(gnd), .Q(regs_12__6_), .vdd(vdd), .CLK(random_clk_bf3__802), .D(_124_), );
  DFFPOSX1 DFFPOSX1_680 (.gnd(gnd), .Q(regs_12__7_), .vdd(vdd), .CLK(random_clk_bf3__1022), .D(_125_), );
  DFFPOSX1 DFFPOSX1_681 (.gnd(gnd), .Q(regs_12__8_), .vdd(vdd), .CLK(random_clk_bf3__1242), .D(_126_), );
  DFFPOSX1 DFFPOSX1_682 (.gnd(gnd), .Q(regs_12__9_), .vdd(vdd), .CLK(random_clk_bf3__1462), .D(_127_), );
  DFFPOSX1 DFFPOSX1_683 (.gnd(gnd), .Q(regs_12__10_), .vdd(vdd), .CLK(random_clk_bf3__1682), .D(_97_), );
  DFFPOSX1 DFFPOSX1_684 (.gnd(gnd), .Q(regs_12__11_), .vdd(vdd), .CLK(random_clk_bf3__1902), .D(_98_), );
  DFFPOSX1 DFFPOSX1_685 (.gnd(gnd), .Q(regs_12__12_), .vdd(vdd), .CLK(random_clk_bf3__182), .D(_99_), );
  DFFPOSX1 DFFPOSX1_686 (.gnd(gnd), .Q(regs_12__13_), .vdd(vdd), .CLK(random_clk_bf3__382), .D(_100_), );
  DFFPOSX1 DFFPOSX1_687 (.gnd(gnd), .Q(regs_12__14_), .vdd(vdd), .CLK(random_clk_bf3__602), .D(_101_), );
  DFFPOSX1 DFFPOSX1_688 (.gnd(gnd), .Q(regs_12__15_), .vdd(vdd), .CLK(random_clk_bf3__822), .D(_102_), );
  DFFPOSX1 DFFPOSX1_689 (.gnd(gnd), .Q(regs_12__16_), .vdd(vdd), .CLK(random_clk_bf3__1042), .D(_103_), );
  DFFPOSX1 DFFPOSX1_690 (.gnd(gnd), .Q(regs_12__17_), .vdd(vdd), .CLK(random_clk_bf3__1262), .D(_104_), );
  DFFPOSX1 DFFPOSX1_691 (.gnd(gnd), .Q(regs_12__18_), .vdd(vdd), .CLK(random_clk_bf3__1482), .D(_105_), );
  DFFPOSX1 DFFPOSX1_692 (.gnd(gnd), .Q(regs_12__19_), .vdd(vdd), .CLK(random_clk_bf3__1702), .D(_106_), );
  DFFPOSX1 DFFPOSX1_693 (.gnd(gnd), .Q(regs_12__20_), .vdd(vdd), .CLK(clock_bf2__28), .D(_108_), );
  DFFPOSX1 DFFPOSX1_694 (.gnd(gnd), .Q(regs_12__21_), .vdd(vdd), .CLK(clock_bf2__7), .D(_109_), );
  DFFPOSX1 DFFPOSX1_695 (.gnd(gnd), .Q(regs_12__22_), .vdd(vdd), .CLK(clock_bf2__18), .D(_110_), );
  DFFPOSX1 DFFPOSX1_696 (.gnd(gnd), .Q(regs_12__23_), .vdd(vdd), .CLK(random_clk_bf3__402), .D(_111_), );
  DFFPOSX1 DFFPOSX1_697 (.gnd(gnd), .Q(regs_12__24_), .vdd(vdd), .CLK(random_clk_bf3__622), .D(_112_), );
  DFFPOSX1 DFFPOSX1_698 (.gnd(gnd), .Q(regs_12__25_), .vdd(vdd), .CLK(random_clk_bf3__842), .D(_113_), );
  DFFPOSX1 DFFPOSX1_699 (.gnd(gnd), .Q(regs_12__26_), .vdd(vdd), .CLK(random_clk_bf3__1062), .D(_114_), );
  DFFPOSX1 DFFPOSX1_700 (.gnd(gnd), .Q(regs_12__27_), .vdd(vdd), .CLK(random_clk_bf3__1282), .D(_115_), );
  DFFPOSX1 DFFPOSX1_701 (.gnd(gnd), .Q(regs_12__28_), .vdd(vdd), .CLK(random_clk_bf3__1502), .D(_116_), );
  DFFPOSX1 DFFPOSX1_702 (.gnd(gnd), .Q(regs_12__29_), .vdd(vdd), .CLK(random_clk_bf3__1722), .D(_117_), );
  DFFPOSX1 DFFPOSX1_703 (.gnd(gnd), .Q(regs_12__30_), .vdd(vdd), .CLK(random_clk_bf3__2), .D(_119_), );
  DFFPOSX1 DFFPOSX1_704 (.gnd(gnd), .Q(regs_12__31_), .vdd(vdd), .CLK(random_clk_bf3__202), .D(_120_), );
  DFFPOSX1 DFFPOSX1_705 (.gnd(gnd), .Q(regs_10__0_), .vdd(vdd), .CLK(random_clk_bf3__422), .D(_32_), );
  DFFPOSX1 DFFPOSX1_706 (.gnd(gnd), .Q(regs_10__1_), .vdd(vdd), .CLK(random_clk_bf3__642), .D(_43_), );
  DFFPOSX1 DFFPOSX1_707 (.gnd(gnd), .Q(regs_10__2_), .vdd(vdd), .CLK(random_clk_bf3__862), .D(_54_), );
  DFFPOSX1 DFFPOSX1_708 (.gnd(gnd), .Q(regs_10__3_), .vdd(vdd), .CLK(random_clk_bf3__1082), .D(_57_), );
  DFFPOSX1 DFFPOSX1_709 (.gnd(gnd), .Q(regs_10__4_), .vdd(vdd), .CLK(random_clk_bf3__1302), .D(_58_), );
  DFFPOSX1 DFFPOSX1_710 (.gnd(gnd), .Q(regs_10__5_), .vdd(vdd), .CLK(random_clk_bf3__1522), .D(_59_), );
  DFFPOSX1 DFFPOSX1_711 (.gnd(gnd), .Q(regs_10__6_), .vdd(vdd), .CLK(random_clk_bf3__1742), .D(_60_), );
  DFFPOSX1 DFFPOSX1_712 (.gnd(gnd), .Q(regs_10__7_), .vdd(vdd), .CLK(random_clk_bf3__22), .D(_61_), );
  DFFPOSX1 DFFPOSX1_713 (.gnd(gnd), .Q(regs_10__8_), .vdd(vdd), .CLK(random_clk_bf3__222), .D(_62_), );
  DFFPOSX1 DFFPOSX1_714 (.gnd(gnd), .Q(regs_10__9_), .vdd(vdd), .CLK(random_clk_bf3__442), .D(_63_), );
  DFFPOSX1 DFFPOSX1_715 (.gnd(gnd), .Q(regs_10__10_), .vdd(vdd), .CLK(random_clk_bf3__662), .D(_33_), );
  DFFPOSX1 DFFPOSX1_716 (.gnd(gnd), .Q(regs_10__11_), .vdd(vdd), .CLK(random_clk_bf3__882), .D(_34_), );
  DFFPOSX1 DFFPOSX1_717 (.gnd(gnd), .Q(regs_10__12_), .vdd(vdd), .CLK(random_clk_bf3__1102), .D(_35_), );
  DFFPOSX1 DFFPOSX1_718 (.gnd(gnd), .Q(regs_10__13_), .vdd(vdd), .CLK(random_clk_bf3__1322), .D(_36_), );
  DFFPOSX1 DFFPOSX1_719 (.gnd(gnd), .Q(regs_10__14_), .vdd(vdd), .CLK(random_clk_bf3__1542), .D(_37_), );
  DFFPOSX1 DFFPOSX1_720 (.gnd(gnd), .Q(regs_10__15_), .vdd(vdd), .CLK(random_clk_bf3__1762), .D(_38_), );
  DFFPOSX1 DFFPOSX1_721 (.gnd(gnd), .Q(regs_10__16_), .vdd(vdd), .CLK(random_clk_bf3__42), .D(_39_), );
  DFFPOSX1 DFFPOSX1_722 (.gnd(gnd), .Q(regs_10__17_), .vdd(vdd), .CLK(random_clk_bf3__242), .D(_40_), );
  DFFPOSX1 DFFPOSX1_723 (.gnd(gnd), .Q(regs_10__18_), .vdd(vdd), .CLK(random_clk_bf3__462), .D(_41_), );
  DFFPOSX1 DFFPOSX1_724 (.gnd(gnd), .Q(regs_10__19_), .vdd(vdd), .CLK(random_clk_bf3__682), .D(_42_), );
  DFFPOSX1 DFFPOSX1_725 (.gnd(gnd), .Q(regs_10__20_), .vdd(vdd), .CLK(random_clk_bf3__902), .D(_44_), );
  DFFPOSX1 DFFPOSX1_726 (.gnd(gnd), .Q(regs_10__21_), .vdd(vdd), .CLK(random_clk_bf3__1122), .D(_45_), );
  DFFPOSX1 DFFPOSX1_727 (.gnd(gnd), .Q(regs_10__22_), .vdd(vdd), .CLK(random_clk_bf3__1342), .D(_46_), );
  DFFPOSX1 DFFPOSX1_728 (.gnd(gnd), .Q(regs_10__23_), .vdd(vdd), .CLK(random_clk_bf3__1562), .D(_47_), );
  DFFPOSX1 DFFPOSX1_729 (.gnd(gnd), .Q(regs_10__24_), .vdd(vdd), .CLK(random_clk_bf3__1782), .D(_48_), );
  DFFPOSX1 DFFPOSX1_730 (.gnd(gnd), .Q(regs_10__25_), .vdd(vdd), .CLK(random_clk_bf3__62), .D(_49_), );
  DFFPOSX1 DFFPOSX1_731 (.gnd(gnd), .Q(regs_10__26_), .vdd(vdd), .CLK(random_clk_bf3__262), .D(_50_), );
  DFFPOSX1 DFFPOSX1_732 (.gnd(gnd), .Q(regs_10__27_), .vdd(vdd), .CLK(random_clk_bf3__482), .D(_51_), );
  DFFPOSX1 DFFPOSX1_733 (.gnd(gnd), .Q(regs_10__28_), .vdd(vdd), .CLK(random_clk_bf3__702), .D(_52_), );
  DFFPOSX1 DFFPOSX1_734 (.gnd(gnd), .Q(regs_10__29_), .vdd(vdd), .CLK(random_clk_bf3__922), .D(_53_), );
  DFFPOSX1 DFFPOSX1_735 (.gnd(gnd), .Q(regs_10__30_), .vdd(vdd), .CLK(random_clk_bf3__1142), .D(_55_), );
  DFFPOSX1 DFFPOSX1_736 (.gnd(gnd), .Q(regs_10__31_), .vdd(vdd), .CLK(random_clk_bf3__1362), .D(_56_), );
  DFFPOSX1 DFFPOSX1_737 (.gnd(gnd), .Q(regs_9__0_), .vdd(vdd), .CLK(random_clk_bf3__1582), .D(_960_), );
  DFFPOSX1 DFFPOSX1_738 (.gnd(gnd), .Q(regs_9__1_), .vdd(vdd), .CLK(random_clk_bf3__1802), .D(_971_), );
  DFFPOSX1 DFFPOSX1_739 (.gnd(gnd), .Q(regs_9__2_), .vdd(vdd), .CLK(random_clk_bf3__82), .D(_982_), );
  DFFPOSX1 DFFPOSX1_740 (.gnd(gnd), .Q(regs_9__3_), .vdd(vdd), .CLK(random_clk_bf3__282), .D(_985_), );
  DFFPOSX1 DFFPOSX1_741 (.gnd(gnd), .Q(regs_9__4_), .vdd(vdd), .CLK(random_clk_bf3__502), .D(_986_), );
  DFFPOSX1 DFFPOSX1_742 (.gnd(gnd), .Q(regs_9__5_), .vdd(vdd), .CLK(random_clk_bf3__722), .D(_987_), );
  DFFPOSX1 DFFPOSX1_743 (.gnd(gnd), .Q(regs_9__6_), .vdd(vdd), .CLK(random_clk_bf3__942), .D(_988_), );
  DFFPOSX1 DFFPOSX1_744 (.gnd(gnd), .Q(regs_9__7_), .vdd(vdd), .CLK(random_clk_bf3__1162), .D(_989_), );
  DFFPOSX1 DFFPOSX1_745 (.gnd(gnd), .Q(regs_9__8_), .vdd(vdd), .CLK(random_clk_bf3__1382), .D(_990_), );
  DFFPOSX1 DFFPOSX1_746 (.gnd(gnd), .Q(regs_9__9_), .vdd(vdd), .CLK(random_clk_bf3__1602), .D(_991_), );
  DFFPOSX1 DFFPOSX1_747 (.gnd(gnd), .Q(regs_9__10_), .vdd(vdd), .CLK(random_clk_bf3__1822), .D(_961_), );
  DFFPOSX1 DFFPOSX1_748 (.gnd(gnd), .Q(regs_9__11_), .vdd(vdd), .CLK(random_clk_bf3__102), .D(_962_), );
  DFFPOSX1 DFFPOSX1_749 (.gnd(gnd), .Q(regs_9__12_), .vdd(vdd), .CLK(random_clk_bf3__302), .D(_963_), );
  DFFPOSX1 DFFPOSX1_750 (.gnd(gnd), .Q(regs_9__13_), .vdd(vdd), .CLK(random_clk_bf3__522), .D(_964_), );
  DFFPOSX1 DFFPOSX1_751 (.gnd(gnd), .Q(regs_9__14_), .vdd(vdd), .CLK(random_clk_bf3__742), .D(_965_), );
  DFFPOSX1 DFFPOSX1_752 (.gnd(gnd), .Q(regs_9__15_), .vdd(vdd), .CLK(random_clk_bf3__962), .D(_966_), );
  DFFPOSX1 DFFPOSX1_753 (.gnd(gnd), .Q(regs_9__16_), .vdd(vdd), .CLK(random_clk_bf3__1182), .D(_967_), );
  DFFPOSX1 DFFPOSX1_754 (.gnd(gnd), .Q(regs_9__17_), .vdd(vdd), .CLK(random_clk_bf3__1402), .D(_968_), );
  DFFPOSX1 DFFPOSX1_755 (.gnd(gnd), .Q(regs_9__18_), .vdd(vdd), .CLK(random_clk_bf3__1622), .D(_969_), );
  DFFPOSX1 DFFPOSX1_756 (.gnd(gnd), .Q(regs_9__19_), .vdd(vdd), .CLK(random_clk_bf3__1842), .D(_970_), );
  DFFPOSX1 DFFPOSX1_757 (.gnd(gnd), .Q(regs_9__20_), .vdd(vdd), .CLK(random_clk_bf3__122), .D(_972_), );
  DFFPOSX1 DFFPOSX1_758 (.gnd(gnd), .Q(regs_9__21_), .vdd(vdd), .CLK(random_clk_bf3__322), .D(_973_), );
  DFFPOSX1 DFFPOSX1_759 (.gnd(gnd), .Q(regs_9__22_), .vdd(vdd), .CLK(random_clk_bf3__542), .D(_974_), );
  DFFPOSX1 DFFPOSX1_760 (.gnd(gnd), .Q(regs_9__23_), .vdd(vdd), .CLK(random_clk_bf3__762), .D(_975_), );
  DFFPOSX1 DFFPOSX1_761 (.gnd(gnd), .Q(regs_9__24_), .vdd(vdd), .CLK(random_clk_bf3__982), .D(_976_), );
  DFFPOSX1 DFFPOSX1_762 (.gnd(gnd), .Q(regs_9__25_), .vdd(vdd), .CLK(random_clk_bf3__1202), .D(_977_), );
  DFFPOSX1 DFFPOSX1_763 (.gnd(gnd), .Q(regs_9__26_), .vdd(vdd), .CLK(random_clk_bf3__1422), .D(_978_), );
  DFFPOSX1 DFFPOSX1_764 (.gnd(gnd), .Q(regs_9__27_), .vdd(vdd), .CLK(random_clk_bf3__1642), .D(_979_), );
  DFFPOSX1 DFFPOSX1_765 (.gnd(gnd), .Q(regs_9__28_), .vdd(vdd), .CLK(random_clk_bf3__1862), .D(_980_), );
  DFFPOSX1 DFFPOSX1_766 (.gnd(gnd), .Q(regs_9__29_), .vdd(vdd), .CLK(random_clk_bf3__142), .D(_981_), );
  DFFPOSX1 DFFPOSX1_767 (.gnd(gnd), .Q(regs_9__30_), .vdd(vdd), .CLK(random_clk_bf3__342), .D(_983_), );
  DFFPOSX1 DFFPOSX1_768 (.gnd(gnd), .Q(regs_9__31_), .vdd(vdd), .CLK(random_clk_bf3__562), .D(_984_), );
  DFFPOSX1 DFFPOSX1_769 (.gnd(gnd), .Q(regs_8__0_), .vdd(vdd), .CLK(random_clk_bf3__782), .D(_928_), );
  DFFPOSX1 DFFPOSX1_770 (.gnd(gnd), .Q(regs_8__1_), .vdd(vdd), .CLK(random_clk_bf3__1002), .D(_939_), );
  DFFPOSX1 DFFPOSX1_771 (.gnd(gnd), .Q(regs_8__2_), .vdd(vdd), .CLK(random_clk_bf3__1222), .D(_950_), );
  DFFPOSX1 DFFPOSX1_772 (.gnd(gnd), .Q(regs_8__3_), .vdd(vdd), .CLK(random_clk_bf3__1442), .D(_953_), );
  DFFPOSX1 DFFPOSX1_773 (.gnd(gnd), .Q(regs_8__4_), .vdd(vdd), .CLK(random_clk_bf3__1662), .D(_954_), );
  DFFPOSX1 DFFPOSX1_774 (.gnd(gnd), .Q(regs_8__5_), .vdd(vdd), .CLK(random_clk_bf3__1882), .D(_955_), );
  DFFPOSX1 DFFPOSX1_775 (.gnd(gnd), .Q(regs_8__6_), .vdd(vdd), .CLK(random_clk_bf3__162), .D(_956_), );
  DFFPOSX1 DFFPOSX1_776 (.gnd(gnd), .Q(regs_8__7_), .vdd(vdd), .CLK(random_clk_bf3__362), .D(_957_), );
  DFFPOSX1 DFFPOSX1_777 (.gnd(gnd), .Q(regs_8__8_), .vdd(vdd), .CLK(random_clk_bf3__582), .D(_958_), );
  DFFPOSX1 DFFPOSX1_778 (.gnd(gnd), .Q(regs_8__9_), .vdd(vdd), .CLK(random_clk_bf3__802), .D(_959_), );
  DFFPOSX1 DFFPOSX1_779 (.gnd(gnd), .Q(regs_8__10_), .vdd(vdd), .CLK(random_clk_bf3__1022), .D(_929_), );
  DFFPOSX1 DFFPOSX1_780 (.gnd(gnd), .Q(regs_8__11_), .vdd(vdd), .CLK(random_clk_bf3__1242), .D(_930_), );
  DFFPOSX1 DFFPOSX1_781 (.gnd(gnd), .Q(regs_8__12_), .vdd(vdd), .CLK(random_clk_bf3__1462), .D(_931_), );
  DFFPOSX1 DFFPOSX1_782 (.gnd(gnd), .Q(regs_8__13_), .vdd(vdd), .CLK(random_clk_bf3__1682), .D(_932_), );
  DFFPOSX1 DFFPOSX1_783 (.gnd(gnd), .Q(regs_8__14_), .vdd(vdd), .CLK(random_clk_bf3__1902), .D(_933_), );
  DFFPOSX1 DFFPOSX1_784 (.gnd(gnd), .Q(regs_8__15_), .vdd(vdd), .CLK(random_clk_bf3__182), .D(_934_), );
  DFFPOSX1 DFFPOSX1_785 (.gnd(gnd), .Q(regs_8__16_), .vdd(vdd), .CLK(random_clk_bf3__382), .D(_935_), );
  DFFPOSX1 DFFPOSX1_786 (.gnd(gnd), .Q(regs_8__17_), .vdd(vdd), .CLK(random_clk_bf3__602), .D(_936_), );
  DFFPOSX1 DFFPOSX1_787 (.gnd(gnd), .Q(regs_8__18_), .vdd(vdd), .CLK(random_clk_bf3__822), .D(_937_), );
  DFFPOSX1 DFFPOSX1_788 (.gnd(gnd), .Q(regs_8__19_), .vdd(vdd), .CLK(random_clk_bf3__1042), .D(_938_), );
  DFFPOSX1 DFFPOSX1_789 (.gnd(gnd), .Q(regs_8__20_), .vdd(vdd), .CLK(random_clk_bf3__1262), .D(_940_), );
  DFFPOSX1 DFFPOSX1_790 (.gnd(gnd), .Q(regs_8__21_), .vdd(vdd), .CLK(random_clk_bf3__1482), .D(_941_), );
  DFFPOSX1 DFFPOSX1_791 (.gnd(gnd), .Q(regs_8__22_), .vdd(vdd), .CLK(random_clk_bf3__1702), .D(_942_), );
  DFFPOSX1 DFFPOSX1_792 (.gnd(gnd), .Q(regs_8__23_), .vdd(vdd), .CLK(clock_bf2__29), .D(_943_), );
  DFFPOSX1 DFFPOSX1_793 (.gnd(gnd), .Q(regs_8__24_), .vdd(vdd), .CLK(clock_bf2__8), .D(_944_), );
  DFFPOSX1 DFFPOSX1_794 (.gnd(gnd), .Q(regs_8__25_), .vdd(vdd), .CLK(clock_bf2__19), .D(_945_), );
  DFFPOSX1 DFFPOSX1_795 (.gnd(gnd), .Q(regs_8__26_), .vdd(vdd), .CLK(random_clk_bf3__402), .D(_946_), );
  DFFPOSX1 DFFPOSX1_796 (.gnd(gnd), .Q(regs_8__27_), .vdd(vdd), .CLK(random_clk_bf3__622), .D(_947_), );
  DFFPOSX1 DFFPOSX1_797 (.gnd(gnd), .Q(regs_8__28_), .vdd(vdd), .CLK(random_clk_bf3__842), .D(_948_), );
  DFFPOSX1 DFFPOSX1_798 (.gnd(gnd), .Q(regs_8__29_), .vdd(vdd), .CLK(random_clk_bf3__1062), .D(_949_), );
  DFFPOSX1 DFFPOSX1_799 (.gnd(gnd), .Q(regs_8__30_), .vdd(vdd), .CLK(random_clk_bf3__1282), .D(_951_), );
  DFFPOSX1 DFFPOSX1_800 (.gnd(gnd), .Q(regs_8__31_), .vdd(vdd), .CLK(random_clk_bf3__1502), .D(_952_), );
  DFFPOSX1 DFFPOSX1_801 (.gnd(gnd), .Q(regs_4__0_), .vdd(vdd), .CLK(random_clk_bf3__1722), .D(_800_), );
  DFFPOSX1 DFFPOSX1_802 (.gnd(gnd), .Q(regs_4__1_), .vdd(vdd), .CLK(random_clk_bf3__2), .D(_811_), );
  DFFPOSX1 DFFPOSX1_803 (.gnd(gnd), .Q(regs_4__2_), .vdd(vdd), .CLK(random_clk_bf3__202), .D(_822_), );
  DFFPOSX1 DFFPOSX1_804 (.gnd(gnd), .Q(regs_4__3_), .vdd(vdd), .CLK(random_clk_bf3__422), .D(_825_), );
  DFFPOSX1 DFFPOSX1_805 (.gnd(gnd), .Q(regs_4__4_), .vdd(vdd), .CLK(random_clk_bf3__642), .D(_826_), );
  DFFPOSX1 DFFPOSX1_806 (.gnd(gnd), .Q(regs_4__5_), .vdd(vdd), .CLK(random_clk_bf3__862), .D(_827_), );
  DFFPOSX1 DFFPOSX1_807 (.gnd(gnd), .Q(regs_4__6_), .vdd(vdd), .CLK(random_clk_bf3__1082), .D(_828_), );
  DFFPOSX1 DFFPOSX1_808 (.gnd(gnd), .Q(regs_4__7_), .vdd(vdd), .CLK(random_clk_bf3__1302), .D(_829_), );
  DFFPOSX1 DFFPOSX1_809 (.gnd(gnd), .Q(regs_4__8_), .vdd(vdd), .CLK(random_clk_bf3__1522), .D(_830_), );
  DFFPOSX1 DFFPOSX1_810 (.gnd(gnd), .Q(regs_4__9_), .vdd(vdd), .CLK(random_clk_bf3__1742), .D(_831_), );
  DFFPOSX1 DFFPOSX1_811 (.gnd(gnd), .Q(regs_4__10_), .vdd(vdd), .CLK(random_clk_bf3__22), .D(_801_), );
  DFFPOSX1 DFFPOSX1_812 (.gnd(gnd), .Q(regs_4__11_), .vdd(vdd), .CLK(random_clk_bf3__222), .D(_802_), );
  DFFPOSX1 DFFPOSX1_813 (.gnd(gnd), .Q(regs_4__12_), .vdd(vdd), .CLK(random_clk_bf3__442), .D(_803_), );
  DFFPOSX1 DFFPOSX1_814 (.gnd(gnd), .Q(regs_4__13_), .vdd(vdd), .CLK(random_clk_bf3__662), .D(_804_), );
  DFFPOSX1 DFFPOSX1_815 (.gnd(gnd), .Q(regs_4__14_), .vdd(vdd), .CLK(random_clk_bf3__882), .D(_805_), );
  DFFPOSX1 DFFPOSX1_816 (.gnd(gnd), .Q(regs_4__15_), .vdd(vdd), .CLK(random_clk_bf3__1102), .D(_806_), );
  DFFPOSX1 DFFPOSX1_817 (.gnd(gnd), .Q(regs_4__16_), .vdd(vdd), .CLK(random_clk_bf3__1322), .D(_807_), );
  DFFPOSX1 DFFPOSX1_818 (.gnd(gnd), .Q(regs_4__17_), .vdd(vdd), .CLK(random_clk_bf3__1542), .D(_808_), );
  DFFPOSX1 DFFPOSX1_819 (.gnd(gnd), .Q(regs_4__18_), .vdd(vdd), .CLK(random_clk_bf3__1762), .D(_809_), );
  DFFPOSX1 DFFPOSX1_820 (.gnd(gnd), .Q(regs_4__19_), .vdd(vdd), .CLK(random_clk_bf3__42), .D(_810_), );
  DFFPOSX1 DFFPOSX1_821 (.gnd(gnd), .Q(regs_4__20_), .vdd(vdd), .CLK(random_clk_bf3__242), .D(_812_), );
  DFFPOSX1 DFFPOSX1_822 (.gnd(gnd), .Q(regs_4__21_), .vdd(vdd), .CLK(random_clk_bf3__462), .D(_813_), );
  DFFPOSX1 DFFPOSX1_823 (.gnd(gnd), .Q(regs_4__22_), .vdd(vdd), .CLK(random_clk_bf3__682), .D(_814_), );
  DFFPOSX1 DFFPOSX1_824 (.gnd(gnd), .Q(regs_4__23_), .vdd(vdd), .CLK(random_clk_bf3__902), .D(_815_), );
  DFFPOSX1 DFFPOSX1_825 (.gnd(gnd), .Q(regs_4__24_), .vdd(vdd), .CLK(random_clk_bf3__1122), .D(_816_), );
  DFFPOSX1 DFFPOSX1_826 (.gnd(gnd), .Q(regs_4__25_), .vdd(vdd), .CLK(random_clk_bf3__1342), .D(_817_), );
  DFFPOSX1 DFFPOSX1_827 (.gnd(gnd), .Q(regs_4__26_), .vdd(vdd), .CLK(random_clk_bf3__1562), .D(_818_), );
  DFFPOSX1 DFFPOSX1_828 (.gnd(gnd), .Q(regs_4__27_), .vdd(vdd), .CLK(random_clk_bf3__1782), .D(_819_), );
  DFFPOSX1 DFFPOSX1_829 (.gnd(gnd), .Q(regs_4__28_), .vdd(vdd), .CLK(random_clk_bf3__62), .D(_820_), );
  DFFPOSX1 DFFPOSX1_830 (.gnd(gnd), .Q(regs_4__29_), .vdd(vdd), .CLK(random_clk_bf3__262), .D(_821_), );
  DFFPOSX1 DFFPOSX1_831 (.gnd(gnd), .Q(regs_4__30_), .vdd(vdd), .CLK(random_clk_bf3__482), .D(_823_), );
  DFFPOSX1 DFFPOSX1_832 (.gnd(gnd), .Q(regs_4__31_), .vdd(vdd), .CLK(random_clk_bf3__702), .D(_824_), );
  DFFPOSX1 DFFPOSX1_833 (.gnd(gnd), .Q(regs_7__0_), .vdd(vdd), .CLK(random_clk_bf3__922), .D(_896_), );
  DFFPOSX1 DFFPOSX1_834 (.gnd(gnd), .Q(regs_7__1_), .vdd(vdd), .CLK(random_clk_bf3__1142), .D(_907_), );
  DFFPOSX1 DFFPOSX1_835 (.gnd(gnd), .Q(regs_7__2_), .vdd(vdd), .CLK(random_clk_bf3__1362), .D(_918_), );
  DFFPOSX1 DFFPOSX1_836 (.gnd(gnd), .Q(regs_7__3_), .vdd(vdd), .CLK(random_clk_bf3__1582), .D(_921_), );
  DFFPOSX1 DFFPOSX1_837 (.gnd(gnd), .Q(regs_7__4_), .vdd(vdd), .CLK(random_clk_bf3__1802), .D(_922_), );
  DFFPOSX1 DFFPOSX1_838 (.gnd(gnd), .Q(regs_7__5_), .vdd(vdd), .CLK(random_clk_bf3__82), .D(_923_), );
  DFFPOSX1 DFFPOSX1_839 (.gnd(gnd), .Q(regs_7__6_), .vdd(vdd), .CLK(random_clk_bf3__282), .D(_924_), );
  DFFPOSX1 DFFPOSX1_840 (.gnd(gnd), .Q(regs_7__7_), .vdd(vdd), .CLK(random_clk_bf3__502), .D(_925_), );
  DFFPOSX1 DFFPOSX1_841 (.gnd(gnd), .Q(regs_7__8_), .vdd(vdd), .CLK(random_clk_bf3__722), .D(_926_), );
  DFFPOSX1 DFFPOSX1_842 (.gnd(gnd), .Q(regs_7__9_), .vdd(vdd), .CLK(random_clk_bf3__942), .D(_927_), );
  DFFPOSX1 DFFPOSX1_843 (.gnd(gnd), .Q(regs_7__10_), .vdd(vdd), .CLK(random_clk_bf3__1162), .D(_897_), );
  DFFPOSX1 DFFPOSX1_844 (.gnd(gnd), .Q(regs_7__11_), .vdd(vdd), .CLK(random_clk_bf3__1382), .D(_898_), );
  DFFPOSX1 DFFPOSX1_845 (.gnd(gnd), .Q(regs_7__12_), .vdd(vdd), .CLK(random_clk_bf3__1602), .D(_899_), );
  DFFPOSX1 DFFPOSX1_846 (.gnd(gnd), .Q(regs_7__13_), .vdd(vdd), .CLK(random_clk_bf3__1822), .D(_900_), );
  DFFPOSX1 DFFPOSX1_847 (.gnd(gnd), .Q(regs_7__14_), .vdd(vdd), .CLK(random_clk_bf3__102), .D(_901_), );
  DFFPOSX1 DFFPOSX1_848 (.gnd(gnd), .Q(regs_7__15_), .vdd(vdd), .CLK(random_clk_bf3__302), .D(_902_), );
  DFFPOSX1 DFFPOSX1_849 (.gnd(gnd), .Q(regs_7__16_), .vdd(vdd), .CLK(random_clk_bf3__522), .D(_903_), );
  DFFPOSX1 DFFPOSX1_850 (.gnd(gnd), .Q(regs_7__17_), .vdd(vdd), .CLK(random_clk_bf3__742), .D(_904_), );
  DFFPOSX1 DFFPOSX1_851 (.gnd(gnd), .Q(regs_7__18_), .vdd(vdd), .CLK(random_clk_bf3__962), .D(_905_), );
  DFFPOSX1 DFFPOSX1_852 (.gnd(gnd), .Q(regs_7__19_), .vdd(vdd), .CLK(random_clk_bf3__1182), .D(_906_), );
  DFFPOSX1 DFFPOSX1_853 (.gnd(gnd), .Q(regs_7__20_), .vdd(vdd), .CLK(random_clk_bf3__1402), .D(_908_), );
  DFFPOSX1 DFFPOSX1_854 (.gnd(gnd), .Q(regs_7__21_), .vdd(vdd), .CLK(random_clk_bf3__1622), .D(_909_), );
  DFFPOSX1 DFFPOSX1_855 (.gnd(gnd), .Q(regs_7__22_), .vdd(vdd), .CLK(random_clk_bf3__1842), .D(_910_), );
  DFFPOSX1 DFFPOSX1_856 (.gnd(gnd), .Q(regs_7__23_), .vdd(vdd), .CLK(random_clk_bf3__122), .D(_911_), );
  DFFPOSX1 DFFPOSX1_857 (.gnd(gnd), .Q(regs_7__24_), .vdd(vdd), .CLK(random_clk_bf3__322), .D(_912_), );
  DFFPOSX1 DFFPOSX1_858 (.gnd(gnd), .Q(regs_7__25_), .vdd(vdd), .CLK(random_clk_bf3__542), .D(_913_), );
  DFFPOSX1 DFFPOSX1_859 (.gnd(gnd), .Q(regs_7__26_), .vdd(vdd), .CLK(random_clk_bf3__762), .D(_914_), );
  DFFPOSX1 DFFPOSX1_860 (.gnd(gnd), .Q(regs_7__27_), .vdd(vdd), .CLK(random_clk_bf3__982), .D(_915_), );
  DFFPOSX1 DFFPOSX1_861 (.gnd(gnd), .Q(regs_7__28_), .vdd(vdd), .CLK(random_clk_bf3__1202), .D(_916_), );
  DFFPOSX1 DFFPOSX1_862 (.gnd(gnd), .Q(regs_7__29_), .vdd(vdd), .CLK(random_clk_bf3__1422), .D(_917_), );
  DFFPOSX1 DFFPOSX1_863 (.gnd(gnd), .Q(regs_7__30_), .vdd(vdd), .CLK(random_clk_bf3__1642), .D(_919_), );
  DFFPOSX1 DFFPOSX1_864 (.gnd(gnd), .Q(regs_7__31_), .vdd(vdd), .CLK(random_clk_bf3__1862), .D(_920_), );
  DFFPOSX1 DFFPOSX1_865 (.gnd(gnd), .Q(regs_3__0_), .vdd(vdd), .CLK(random_clk_bf3__142), .D(_768_), );
  DFFPOSX1 DFFPOSX1_866 (.gnd(gnd), .Q(regs_3__1_), .vdd(vdd), .CLK(random_clk_bf3__342), .D(_779_), );
  DFFPOSX1 DFFPOSX1_867 (.gnd(gnd), .Q(regs_3__2_), .vdd(vdd), .CLK(random_clk_bf3__562), .D(_790_), );
  DFFPOSX1 DFFPOSX1_868 (.gnd(gnd), .Q(regs_3__3_), .vdd(vdd), .CLK(random_clk_bf3__782), .D(_793_), );
  DFFPOSX1 DFFPOSX1_869 (.gnd(gnd), .Q(regs_3__4_), .vdd(vdd), .CLK(random_clk_bf3__1002), .D(_794_), );
  DFFPOSX1 DFFPOSX1_870 (.gnd(gnd), .Q(regs_3__5_), .vdd(vdd), .CLK(random_clk_bf3__1222), .D(_795_), );
  DFFPOSX1 DFFPOSX1_871 (.gnd(gnd), .Q(regs_3__6_), .vdd(vdd), .CLK(random_clk_bf3__1442), .D(_796_), );
  DFFPOSX1 DFFPOSX1_872 (.gnd(gnd), .Q(regs_3__7_), .vdd(vdd), .CLK(random_clk_bf3__1662), .D(_797_), );
  DFFPOSX1 DFFPOSX1_873 (.gnd(gnd), .Q(regs_3__8_), .vdd(vdd), .CLK(random_clk_bf3__1882), .D(_798_), );
  DFFPOSX1 DFFPOSX1_874 (.gnd(gnd), .Q(regs_3__9_), .vdd(vdd), .CLK(random_clk_bf3__162), .D(_799_), );
  DFFPOSX1 DFFPOSX1_875 (.gnd(gnd), .Q(regs_3__10_), .vdd(vdd), .CLK(random_clk_bf3__362), .D(_769_), );
  DFFPOSX1 DFFPOSX1_876 (.gnd(gnd), .Q(regs_3__11_), .vdd(vdd), .CLK(random_clk_bf3__582), .D(_770_), );
  DFFPOSX1 DFFPOSX1_877 (.gnd(gnd), .Q(regs_3__12_), .vdd(vdd), .CLK(random_clk_bf3__802), .D(_771_), );
  DFFPOSX1 DFFPOSX1_878 (.gnd(gnd), .Q(regs_3__13_), .vdd(vdd), .CLK(random_clk_bf3__1022), .D(_772_), );
  DFFPOSX1 DFFPOSX1_879 (.gnd(gnd), .Q(regs_3__14_), .vdd(vdd), .CLK(random_clk_bf3__1242), .D(_773_), );
  DFFPOSX1 DFFPOSX1_880 (.gnd(gnd), .Q(regs_3__15_), .vdd(vdd), .CLK(random_clk_bf3__1462), .D(_774_), );
  DFFPOSX1 DFFPOSX1_881 (.gnd(gnd), .Q(regs_3__16_), .vdd(vdd), .CLK(random_clk_bf3__1682), .D(_775_), );
  DFFPOSX1 DFFPOSX1_882 (.gnd(gnd), .Q(regs_3__17_), .vdd(vdd), .CLK(random_clk_bf3__1902), .D(_776_), );
  DFFPOSX1 DFFPOSX1_883 (.gnd(gnd), .Q(regs_3__18_), .vdd(vdd), .CLK(random_clk_bf3__182), .D(_777_), );
  DFFPOSX1 DFFPOSX1_884 (.gnd(gnd), .Q(regs_3__19_), .vdd(vdd), .CLK(random_clk_bf3__382), .D(_778_), );
  DFFPOSX1 DFFPOSX1_885 (.gnd(gnd), .Q(regs_3__20_), .vdd(vdd), .CLK(random_clk_bf3__602), .D(_780_), );
  DFFPOSX1 DFFPOSX1_886 (.gnd(gnd), .Q(regs_3__21_), .vdd(vdd), .CLK(random_clk_bf3__822), .D(_781_), );
  DFFPOSX1 DFFPOSX1_887 (.gnd(gnd), .Q(regs_3__22_), .vdd(vdd), .CLK(random_clk_bf3__1042), .D(_782_), );
  DFFPOSX1 DFFPOSX1_888 (.gnd(gnd), .Q(regs_3__23_), .vdd(vdd), .CLK(random_clk_bf3__1262), .D(_783_), );
  DFFPOSX1 DFFPOSX1_889 (.gnd(gnd), .Q(regs_3__24_), .vdd(vdd), .CLK(random_clk_bf3__1482), .D(_784_), );
  DFFPOSX1 DFFPOSX1_890 (.gnd(gnd), .Q(regs_3__25_), .vdd(vdd), .CLK(random_clk_bf3__1702), .D(_785_), );
  DFFPOSX1 DFFPOSX1_891 (.gnd(gnd), .Q(regs_3__26_), .vdd(vdd), .CLK(clock_bf2__30), .D(_786_), );
  DFFPOSX1 DFFPOSX1_892 (.gnd(gnd), .Q(regs_3__27_), .vdd(vdd), .CLK(clock_bf2__9), .D(_787_), );
  DFFPOSX1 DFFPOSX1_893 (.gnd(gnd), .Q(regs_3__28_), .vdd(vdd), .CLK(clock_bf2__20), .D(_788_), );
  DFFPOSX1 DFFPOSX1_894 (.gnd(gnd), .Q(regs_3__29_), .vdd(vdd), .CLK(random_clk_bf3__402), .D(_789_), );
  DFFPOSX1 DFFPOSX1_895 (.gnd(gnd), .Q(regs_3__30_), .vdd(vdd), .CLK(random_clk_bf3__622), .D(_791_), );
  DFFPOSX1 DFFPOSX1_896 (.gnd(gnd), .Q(regs_3__31_), .vdd(vdd), .CLK(random_clk_bf3__842), .D(_792_), );
  DFFPOSX1 DFFPOSX1_897 (.gnd(gnd), .Q(regs_2__0_), .vdd(vdd), .CLK(random_clk_bf3__1062), .D(_704_), );
  DFFPOSX1 DFFPOSX1_898 (.gnd(gnd), .Q(regs_2__1_), .vdd(vdd), .CLK(random_clk_bf3__1282), .D(_715_), );
  DFFPOSX1 DFFPOSX1_899 (.gnd(gnd), .Q(regs_2__2_), .vdd(vdd), .CLK(random_clk_bf3__1502), .D(_726_), );
  DFFPOSX1 DFFPOSX1_900 (.gnd(gnd), .Q(regs_2__3_), .vdd(vdd), .CLK(random_clk_bf3__1722), .D(_729_), );
  DFFPOSX1 DFFPOSX1_901 (.gnd(gnd), .Q(regs_2__4_), .vdd(vdd), .CLK(random_clk_bf3__2), .D(_730_), );
  DFFPOSX1 DFFPOSX1_902 (.gnd(gnd), .Q(regs_2__5_), .vdd(vdd), .CLK(random_clk_bf3__202), .D(_731_), );
  DFFPOSX1 DFFPOSX1_903 (.gnd(gnd), .Q(regs_2__6_), .vdd(vdd), .CLK(random_clk_bf3__422), .D(_732_), );
  DFFPOSX1 DFFPOSX1_904 (.gnd(gnd), .Q(regs_2__7_), .vdd(vdd), .CLK(random_clk_bf3__642), .D(_733_), );
  DFFPOSX1 DFFPOSX1_905 (.gnd(gnd), .Q(regs_2__8_), .vdd(vdd), .CLK(random_clk_bf3__862), .D(_734_), );
  DFFPOSX1 DFFPOSX1_906 (.gnd(gnd), .Q(regs_2__9_), .vdd(vdd), .CLK(random_clk_bf3__1082), .D(_735_), );
  DFFPOSX1 DFFPOSX1_907 (.gnd(gnd), .Q(regs_2__10_), .vdd(vdd), .CLK(random_clk_bf3__1302), .D(_705_), );
  DFFPOSX1 DFFPOSX1_908 (.gnd(gnd), .Q(regs_2__11_), .vdd(vdd), .CLK(random_clk_bf3__1522), .D(_706_), );
  DFFPOSX1 DFFPOSX1_909 (.gnd(gnd), .Q(regs_2__12_), .vdd(vdd), .CLK(random_clk_bf3__1742), .D(_707_), );
  DFFPOSX1 DFFPOSX1_910 (.gnd(gnd), .Q(regs_2__13_), .vdd(vdd), .CLK(random_clk_bf3__22), .D(_708_), );
  DFFPOSX1 DFFPOSX1_911 (.gnd(gnd), .Q(regs_2__14_), .vdd(vdd), .CLK(random_clk_bf3__222), .D(_709_), );
  DFFPOSX1 DFFPOSX1_912 (.gnd(gnd), .Q(regs_2__15_), .vdd(vdd), .CLK(random_clk_bf3__442), .D(_710_), );
  DFFPOSX1 DFFPOSX1_913 (.gnd(gnd), .Q(regs_2__16_), .vdd(vdd), .CLK(random_clk_bf3__662), .D(_711_), );
  DFFPOSX1 DFFPOSX1_914 (.gnd(gnd), .Q(regs_2__17_), .vdd(vdd), .CLK(random_clk_bf3__882), .D(_712_), );
  DFFPOSX1 DFFPOSX1_915 (.gnd(gnd), .Q(regs_2__18_), .vdd(vdd), .CLK(random_clk_bf3__1102), .D(_713_), );
  DFFPOSX1 DFFPOSX1_916 (.gnd(gnd), .Q(regs_2__19_), .vdd(vdd), .CLK(random_clk_bf3__1322), .D(_714_), );
  DFFPOSX1 DFFPOSX1_917 (.gnd(gnd), .Q(regs_2__20_), .vdd(vdd), .CLK(random_clk_bf3__1542), .D(_716_), );
  DFFPOSX1 DFFPOSX1_918 (.gnd(gnd), .Q(regs_2__21_), .vdd(vdd), .CLK(random_clk_bf3__1762), .D(_717_), );
  DFFPOSX1 DFFPOSX1_919 (.gnd(gnd), .Q(regs_2__22_), .vdd(vdd), .CLK(random_clk_bf3__42), .D(_718_), );
  DFFPOSX1 DFFPOSX1_920 (.gnd(gnd), .Q(regs_2__23_), .vdd(vdd), .CLK(random_clk_bf3__242), .D(_719_), );
  DFFPOSX1 DFFPOSX1_921 (.gnd(gnd), .Q(regs_2__24_), .vdd(vdd), .CLK(random_clk_bf3__462), .D(_720_), );
  DFFPOSX1 DFFPOSX1_922 (.gnd(gnd), .Q(regs_2__25_), .vdd(vdd), .CLK(random_clk_bf3__682), .D(_721_), );
  DFFPOSX1 DFFPOSX1_923 (.gnd(gnd), .Q(regs_2__26_), .vdd(vdd), .CLK(random_clk_bf3__902), .D(_722_), );
  DFFPOSX1 DFFPOSX1_924 (.gnd(gnd), .Q(regs_2__27_), .vdd(vdd), .CLK(random_clk_bf3__1122), .D(_723_), );
  DFFPOSX1 DFFPOSX1_925 (.gnd(gnd), .Q(regs_2__28_), .vdd(vdd), .CLK(random_clk_bf3__1342), .D(_724_), );
  DFFPOSX1 DFFPOSX1_926 (.gnd(gnd), .Q(regs_2__29_), .vdd(vdd), .CLK(random_clk_bf3__1562), .D(_725_), );
  DFFPOSX1 DFFPOSX1_927 (.gnd(gnd), .Q(regs_2__30_), .vdd(vdd), .CLK(random_clk_bf3__1782), .D(_727_), );
  DFFPOSX1 DFFPOSX1_928 (.gnd(gnd), .Q(regs_2__31_), .vdd(vdd), .CLK(random_clk_bf3__62), .D(_728_), );
  DFFPOSX1 DFFPOSX1_929 (.gnd(gnd), .Q(regs_6__0_), .vdd(vdd), .CLK(random_clk_bf3__262), .D(_864_), );
  DFFPOSX1 DFFPOSX1_930 (.gnd(gnd), .Q(regs_6__1_), .vdd(vdd), .CLK(random_clk_bf3__482), .D(_875_), );
  DFFPOSX1 DFFPOSX1_931 (.gnd(gnd), .Q(regs_6__2_), .vdd(vdd), .CLK(random_clk_bf3__702), .D(_886_), );
  DFFPOSX1 DFFPOSX1_932 (.gnd(gnd), .Q(regs_6__3_), .vdd(vdd), .CLK(random_clk_bf3__922), .D(_889_), );
  DFFPOSX1 DFFPOSX1_933 (.gnd(gnd), .Q(regs_6__4_), .vdd(vdd), .CLK(random_clk_bf3__1142), .D(_890_), );
  DFFPOSX1 DFFPOSX1_934 (.gnd(gnd), .Q(regs_6__5_), .vdd(vdd), .CLK(random_clk_bf3__1362), .D(_891_), );
  DFFPOSX1 DFFPOSX1_935 (.gnd(gnd), .Q(regs_6__6_), .vdd(vdd), .CLK(random_clk_bf3__1582), .D(_892_), );
  DFFPOSX1 DFFPOSX1_936 (.gnd(gnd), .Q(regs_6__7_), .vdd(vdd), .CLK(random_clk_bf3__1802), .D(_893_), );
  DFFPOSX1 DFFPOSX1_937 (.gnd(gnd), .Q(regs_6__8_), .vdd(vdd), .CLK(random_clk_bf3__82), .D(_894_), );
  DFFPOSX1 DFFPOSX1_938 (.gnd(gnd), .Q(regs_6__9_), .vdd(vdd), .CLK(random_clk_bf3__282), .D(_895_), );
  DFFPOSX1 DFFPOSX1_939 (.gnd(gnd), .Q(regs_6__10_), .vdd(vdd), .CLK(random_clk_bf3__502), .D(_865_), );
  DFFPOSX1 DFFPOSX1_940 (.gnd(gnd), .Q(regs_6__11_), .vdd(vdd), .CLK(random_clk_bf3__722), .D(_866_), );
  DFFPOSX1 DFFPOSX1_941 (.gnd(gnd), .Q(regs_6__12_), .vdd(vdd), .CLK(random_clk_bf3__942), .D(_867_), );
  DFFPOSX1 DFFPOSX1_942 (.gnd(gnd), .Q(regs_6__13_), .vdd(vdd), .CLK(random_clk_bf3__1162), .D(_868_), );
  DFFPOSX1 DFFPOSX1_943 (.gnd(gnd), .Q(regs_6__14_), .vdd(vdd), .CLK(random_clk_bf3__1382), .D(_869_), );
  DFFPOSX1 DFFPOSX1_944 (.gnd(gnd), .Q(regs_6__15_), .vdd(vdd), .CLK(random_clk_bf3__1602), .D(_870_), );
  DFFPOSX1 DFFPOSX1_945 (.gnd(gnd), .Q(regs_6__16_), .vdd(vdd), .CLK(random_clk_bf3__1822), .D(_871_), );
  DFFPOSX1 DFFPOSX1_946 (.gnd(gnd), .Q(regs_6__17_), .vdd(vdd), .CLK(random_clk_bf3__102), .D(_872_), );
  DFFPOSX1 DFFPOSX1_947 (.gnd(gnd), .Q(regs_6__18_), .vdd(vdd), .CLK(random_clk_bf3__302), .D(_873_), );
  DFFPOSX1 DFFPOSX1_948 (.gnd(gnd), .Q(regs_6__19_), .vdd(vdd), .CLK(random_clk_bf3__522), .D(_874_), );
  DFFPOSX1 DFFPOSX1_949 (.gnd(gnd), .Q(regs_6__20_), .vdd(vdd), .CLK(random_clk_bf3__742), .D(_876_), );
  DFFPOSX1 DFFPOSX1_950 (.gnd(gnd), .Q(regs_6__21_), .vdd(vdd), .CLK(random_clk_bf3__962), .D(_877_), );
  DFFPOSX1 DFFPOSX1_951 (.gnd(gnd), .Q(regs_6__22_), .vdd(vdd), .CLK(random_clk_bf3__1182), .D(_878_), );
  DFFPOSX1 DFFPOSX1_952 (.gnd(gnd), .Q(regs_6__23_), .vdd(vdd), .CLK(random_clk_bf3__1402), .D(_879_), );
  DFFPOSX1 DFFPOSX1_953 (.gnd(gnd), .Q(regs_6__24_), .vdd(vdd), .CLK(random_clk_bf3__1622), .D(_880_), );
  DFFPOSX1 DFFPOSX1_954 (.gnd(gnd), .Q(regs_6__25_), .vdd(vdd), .CLK(random_clk_bf3__1842), .D(_881_), );
  DFFPOSX1 DFFPOSX1_955 (.gnd(gnd), .Q(regs_6__26_), .vdd(vdd), .CLK(random_clk_bf3__122), .D(_882_), );
  DFFPOSX1 DFFPOSX1_956 (.gnd(gnd), .Q(regs_6__27_), .vdd(vdd), .CLK(random_clk_bf3__322), .D(_883_), );
  DFFPOSX1 DFFPOSX1_957 (.gnd(gnd), .Q(regs_6__28_), .vdd(vdd), .CLK(random_clk_bf3__542), .D(_884_), );
  DFFPOSX1 DFFPOSX1_958 (.gnd(gnd), .Q(regs_6__29_), .vdd(vdd), .CLK(random_clk_bf3__762), .D(_885_), );
  DFFPOSX1 DFFPOSX1_959 (.gnd(gnd), .Q(regs_6__30_), .vdd(vdd), .CLK(random_clk_bf3__982), .D(_887_), );
  DFFPOSX1 DFFPOSX1_960 (.gnd(gnd), .Q(regs_6__31_), .vdd(vdd), .CLK(random_clk_bf3__1202), .D(_888_), );
  DFFPOSX1 DFFPOSX1_961 (.gnd(gnd), .Q(regs_5__0_), .vdd(vdd), .CLK(random_clk_bf3__1422), .D(_832_), );
  DFFPOSX1 DFFPOSX1_962 (.gnd(gnd), .Q(regs_5__1_), .vdd(vdd), .CLK(random_clk_bf3__1642), .D(_843_), );
  DFFPOSX1 DFFPOSX1_963 (.gnd(gnd), .Q(regs_5__2_), .vdd(vdd), .CLK(random_clk_bf3__1862), .D(_854_), );
  DFFPOSX1 DFFPOSX1_964 (.gnd(gnd), .Q(regs_5__3_), .vdd(vdd), .CLK(random_clk_bf3__142), .D(_857_), );
  DFFPOSX1 DFFPOSX1_965 (.gnd(gnd), .Q(regs_5__4_), .vdd(vdd), .CLK(random_clk_bf3__342), .D(_858_), );
  DFFPOSX1 DFFPOSX1_966 (.gnd(gnd), .Q(regs_5__5_), .vdd(vdd), .CLK(random_clk_bf3__562), .D(_859_), );
  DFFPOSX1 DFFPOSX1_967 (.gnd(gnd), .Q(regs_5__6_), .vdd(vdd), .CLK(random_clk_bf3__782), .D(_860_), );
  DFFPOSX1 DFFPOSX1_968 (.gnd(gnd), .Q(regs_5__7_), .vdd(vdd), .CLK(random_clk_bf3__1002), .D(_861_), );
  DFFPOSX1 DFFPOSX1_969 (.gnd(gnd), .Q(regs_5__8_), .vdd(vdd), .CLK(random_clk_bf3__1222), .D(_862_), );
  DFFPOSX1 DFFPOSX1_970 (.gnd(gnd), .Q(regs_5__9_), .vdd(vdd), .CLK(random_clk_bf3__1442), .D(_863_), );
  DFFPOSX1 DFFPOSX1_971 (.gnd(gnd), .Q(regs_5__10_), .vdd(vdd), .CLK(random_clk_bf3__1662), .D(_833_), );
  DFFPOSX1 DFFPOSX1_972 (.gnd(gnd), .Q(regs_5__11_), .vdd(vdd), .CLK(random_clk_bf3__1882), .D(_834_), );
  DFFPOSX1 DFFPOSX1_973 (.gnd(gnd), .Q(regs_5__12_), .vdd(vdd), .CLK(random_clk_bf3__162), .D(_835_), );
  DFFPOSX1 DFFPOSX1_974 (.gnd(gnd), .Q(regs_5__13_), .vdd(vdd), .CLK(random_clk_bf3__362), .D(_836_), );
  DFFPOSX1 DFFPOSX1_975 (.gnd(gnd), .Q(regs_5__14_), .vdd(vdd), .CLK(random_clk_bf3__582), .D(_837_), );
  DFFPOSX1 DFFPOSX1_976 (.gnd(gnd), .Q(regs_5__15_), .vdd(vdd), .CLK(random_clk_bf3__802), .D(_838_), );
  DFFPOSX1 DFFPOSX1_977 (.gnd(gnd), .Q(regs_5__16_), .vdd(vdd), .CLK(random_clk_bf3__1022), .D(_839_), );
  DFFPOSX1 DFFPOSX1_978 (.gnd(gnd), .Q(regs_5__17_), .vdd(vdd), .CLK(random_clk_bf3__1242), .D(_840_), );
  DFFPOSX1 DFFPOSX1_979 (.gnd(gnd), .Q(regs_5__18_), .vdd(vdd), .CLK(random_clk_bf3__1462), .D(_841_), );
  DFFPOSX1 DFFPOSX1_980 (.gnd(gnd), .Q(regs_5__19_), .vdd(vdd), .CLK(random_clk_bf3__1682), .D(_842_), );
  DFFPOSX1 DFFPOSX1_981 (.gnd(gnd), .Q(regs_5__20_), .vdd(vdd), .CLK(random_clk_bf3__1902), .D(_844_), );
  DFFPOSX1 DFFPOSX1_982 (.gnd(gnd), .Q(regs_5__21_), .vdd(vdd), .CLK(random_clk_bf3__182), .D(_845_), );
  DFFPOSX1 DFFPOSX1_983 (.gnd(gnd), .Q(regs_5__22_), .vdd(vdd), .CLK(random_clk_bf3__382), .D(_846_), );
  DFFPOSX1 DFFPOSX1_984 (.gnd(gnd), .Q(regs_5__23_), .vdd(vdd), .CLK(random_clk_bf3__602), .D(_847_), );
  DFFPOSX1 DFFPOSX1_985 (.gnd(gnd), .Q(regs_5__24_), .vdd(vdd), .CLK(random_clk_bf3__822), .D(_848_), );
  DFFPOSX1 DFFPOSX1_986 (.gnd(gnd), .Q(regs_5__25_), .vdd(vdd), .CLK(random_clk_bf3__1042), .D(_849_), );
  DFFPOSX1 DFFPOSX1_987 (.gnd(gnd), .Q(regs_5__26_), .vdd(vdd), .CLK(random_clk_bf3__1262), .D(_850_), );
  DFFPOSX1 DFFPOSX1_988 (.gnd(gnd), .Q(regs_5__27_), .vdd(vdd), .CLK(random_clk_bf3__1482), .D(_851_), );
  DFFPOSX1 DFFPOSX1_989 (.gnd(gnd), .Q(regs_5__28_), .vdd(vdd), .CLK(random_clk_bf3__1702), .D(_852_), );
  DFFPOSX1 DFFPOSX1_990 (.gnd(gnd), .Q(regs_5__29_), .vdd(vdd), .CLK(clock_bf2__31), .D(_853_), );
  DFFPOSX1 DFFPOSX1_991 (.gnd(gnd), .Q(regs_5__30_), .vdd(vdd), .CLK(clock_bf2__10), .D(_855_), );
  DFFPOSX1 DFFPOSX1_992 (.gnd(gnd), .Q(regs_5__31_), .vdd(vdd), .CLK(clock_bf2__21), .D(_856_), );
  OAI21X1 OAI21X1_458 (.gnd(gnd), .A(_1936_), .Y(_72_), .vdd(vdd), .B(_1902__bF_buf4), .C(_1937_), );
  INVX2 INVX2_211 (.gnd(gnd), .A(regs_11__18_), .Y(_1938_), .vdd(vdd), );
  NAND2X1 NAND2X1_213 (.gnd(gnd), .A(wdata[18]), .Y(_1939_), .vdd(vdd), .B(_1902__bF_buf3), );
  OAI21X1 OAI21X1_459 (.gnd(gnd), .A(_1938_), .Y(_73_), .vdd(vdd), .B(_1902__bF_buf2), .C(_1939_), );
  INVX2 INVX2_212 (.gnd(gnd), .A(regs_11__19_), .Y(_1940_), .vdd(vdd), );
  NAND2X1 NAND2X1_214 (.gnd(gnd), .A(wdata[19]), .Y(_1941_), .vdd(vdd), .B(_1902__bF_buf1), );
  OAI21X1 OAI21X1_460 (.gnd(gnd), .A(_1940_), .Y(_74_), .vdd(vdd), .B(_1902__bF_buf0), .C(_1941_), );
  INVX2 INVX2_213 (.gnd(gnd), .A(regs_11__20_), .Y(_1942_), .vdd(vdd), );
  NAND2X1 NAND2X1_215 (.gnd(gnd), .A(wdata[20]), .Y(_1943_), .vdd(vdd), .B(_1902__bF_buf7), );
  OAI21X1 OAI21X1_461 (.gnd(gnd), .A(_1942_), .Y(_76_), .vdd(vdd), .B(_1902__bF_buf6), .C(_1943_), );
  INVX2 INVX2_214 (.gnd(gnd), .A(regs_11__21_), .Y(_1944_), .vdd(vdd), );
  NAND2X1 NAND2X1_216 (.gnd(gnd), .A(wdata[21]), .Y(_1945_), .vdd(vdd), .B(_1902__bF_buf5), );
  OAI21X1 OAI21X1_462 (.gnd(gnd), .A(_1944_), .Y(_77_), .vdd(vdd), .B(_1902__bF_buf4), .C(_1945_), );
  INVX2 INVX2_215 (.gnd(gnd), .A(regs_11__22_), .Y(_1946_), .vdd(vdd), );
  NAND2X1 NAND2X1_217 (.gnd(gnd), .A(wdata[22]), .Y(_1947_), .vdd(vdd), .B(_1902__bF_buf3), );
  OAI21X1 OAI21X1_463 (.gnd(gnd), .A(_1946_), .Y(_78_), .vdd(vdd), .B(_1902__bF_buf2), .C(_1947_), );
  INVX2 INVX2_216 (.gnd(gnd), .A(regs_11__23_), .Y(_1948_), .vdd(vdd), );
  NAND2X1 NAND2X1_218 (.gnd(gnd), .A(wdata[23]), .Y(_1949_), .vdd(vdd), .B(_1902__bF_buf1), );
  OAI21X1 OAI21X1_464 (.gnd(gnd), .A(_1948_), .Y(_79_), .vdd(vdd), .B(_1902__bF_buf0), .C(_1949_), );
  INVX2 INVX2_217 (.gnd(gnd), .A(regs_11__24_), .Y(_1950_), .vdd(vdd), );
  NAND2X1 NAND2X1_219 (.gnd(gnd), .A(wdata[24]), .Y(_1951_), .vdd(vdd), .B(_1902__bF_buf7), );
  OAI21X1 OAI21X1_465 (.gnd(gnd), .A(_1950_), .Y(_80_), .vdd(vdd), .B(_1902__bF_buf6), .C(_1951_), );
  INVX2 INVX2_218 (.gnd(gnd), .A(regs_11__25_), .Y(_1952_), .vdd(vdd), );
  NAND2X1 NAND2X1_220 (.gnd(gnd), .A(wdata[25]), .Y(_1953_), .vdd(vdd), .B(_1902__bF_buf5), );
  OAI21X1 OAI21X1_466 (.gnd(gnd), .A(_1952_), .Y(_81_), .vdd(vdd), .B(_1902__bF_buf4), .C(_1953_), );
  INVX2 INVX2_219 (.gnd(gnd), .A(regs_11__26_), .Y(_1954_), .vdd(vdd), );
  NAND2X1 NAND2X1_221 (.gnd(gnd), .A(wdata[26]), .Y(_1955_), .vdd(vdd), .B(_1902__bF_buf3), );
  OAI21X1 OAI21X1_467 (.gnd(gnd), .A(_1954_), .Y(_82_), .vdd(vdd), .B(_1902__bF_buf2), .C(_1955_), );
  INVX2 INVX2_220 (.gnd(gnd), .A(regs_11__27_), .Y(_1956_), .vdd(vdd), );
  NAND2X1 NAND2X1_222 (.gnd(gnd), .A(wdata[27]), .Y(_1957_), .vdd(vdd), .B(_1902__bF_buf1), );
  OAI21X1 OAI21X1_468 (.gnd(gnd), .A(_1956_), .Y(_83_), .vdd(vdd), .B(_1902__bF_buf0), .C(_1957_), );
  INVX2 INVX2_221 (.gnd(gnd), .A(regs_11__28_), .Y(_1958_), .vdd(vdd), );
  NAND2X1 NAND2X1_223 (.gnd(gnd), .A(wdata[28]), .Y(_1959_), .vdd(vdd), .B(_1902__bF_buf7), );
  OAI21X1 OAI21X1_469 (.gnd(gnd), .A(_1958_), .Y(_84_), .vdd(vdd), .B(_1902__bF_buf6), .C(_1959_), );
  INVX2 INVX2_222 (.gnd(gnd), .A(regs_11__29_), .Y(_1960_), .vdd(vdd), );
  NAND2X1 NAND2X1_224 (.gnd(gnd), .A(wdata[29]), .Y(_1961_), .vdd(vdd), .B(_1902__bF_buf5), );
  OAI21X1 OAI21X1_470 (.gnd(gnd), .A(_1960_), .Y(_85_), .vdd(vdd), .B(_1902__bF_buf4), .C(_1961_), );
  INVX2 INVX2_223 (.gnd(gnd), .A(regs_11__30_), .Y(_1962_), .vdd(vdd), );
  NAND2X1 NAND2X1_225 (.gnd(gnd), .A(wdata[30]), .Y(_1963_), .vdd(vdd), .B(_1902__bF_buf3), );
  OAI21X1 OAI21X1_471 (.gnd(gnd), .A(_1962_), .Y(_87_), .vdd(vdd), .B(_1902__bF_buf2), .C(_1963_), );
  INVX2 INVX2_224 (.gnd(gnd), .A(regs_11__31_), .Y(_1964_), .vdd(vdd), );
  NAND2X1 NAND2X1_226 (.gnd(gnd), .A(wdata[31]), .Y(_1965_), .vdd(vdd), .B(_1902__bF_buf1), );
  OAI21X1 OAI21X1_472 (.gnd(gnd), .A(_1964_), .Y(_88_), .vdd(vdd), .B(_1902__bF_buf0), .C(_1965_), );
  NOR2X1 NOR2X1_107 (.gnd(gnd), .A(_1001__bF_buf6), .Y(_1966_), .vdd(vdd), .B(_1901__bF_buf4), );
  NOR2X1 NOR2X1_108 (.gnd(gnd), .A(regs_10__0_), .Y(_1967_), .vdd(vdd), .B(_1966__bF_buf7), );
  AOI21X1 AOI21X1_97 (.gnd(gnd), .A(_992__bF_buf1), .Y(_32_), .vdd(vdd), .B(_1966__bF_buf6), .C(_1967_), );
  NOR2X1 NOR2X1_109 (.gnd(gnd), .A(regs_10__1_), .Y(_1968_), .vdd(vdd), .B(_1966__bF_buf5), );
  AOI21X1 AOI21X1_98 (.gnd(gnd), .A(_1003__bF_buf1), .Y(_43_), .vdd(vdd), .B(_1966__bF_buf4), .C(_1968_), );
  NOR2X1 NOR2X1_110 (.gnd(gnd), .A(regs_10__2_), .Y(_1969_), .vdd(vdd), .B(_1966__bF_buf3), );
  AOI21X1 AOI21X1_99 (.gnd(gnd), .A(_1005__bF_buf1), .Y(_54_), .vdd(vdd), .B(_1966__bF_buf2), .C(_1969_), );
  NOR2X1 NOR2X1_111 (.gnd(gnd), .A(regs_10__3_), .Y(_1970_), .vdd(vdd), .B(_1966__bF_buf1), );
  AOI21X1 AOI21X1_100 (.gnd(gnd), .A(_1007__bF_buf1), .Y(_57_), .vdd(vdd), .B(_1966__bF_buf0), .C(_1970_), );
  NOR2X1 NOR2X1_112 (.gnd(gnd), .A(regs_10__4_), .Y(_1971_), .vdd(vdd), .B(_1966__bF_buf7), );
  AOI21X1 AOI21X1_101 (.gnd(gnd), .A(_1009__bF_buf0), .Y(_58_), .vdd(vdd), .B(_1966__bF_buf6), .C(_1971_), );
  NOR2X1 NOR2X1_113 (.gnd(gnd), .A(regs_10__5_), .Y(_1972_), .vdd(vdd), .B(_1966__bF_buf5), );
  AOI21X1 AOI21X1_102 (.gnd(gnd), .A(_1011__bF_buf0), .Y(_59_), .vdd(vdd), .B(_1966__bF_buf4), .C(_1972_), );
  NOR2X1 NOR2X1_114 (.gnd(gnd), .A(regs_10__6_), .Y(_1973_), .vdd(vdd), .B(_1966__bF_buf3), );
  AOI21X1 AOI21X1_103 (.gnd(gnd), .A(_1013__bF_buf0), .Y(_60_), .vdd(vdd), .B(_1966__bF_buf2), .C(_1973_), );
  NOR2X1 NOR2X1_115 (.gnd(gnd), .A(regs_10__7_), .Y(_1974_), .vdd(vdd), .B(_1966__bF_buf1), );
  AOI21X1 AOI21X1_104 (.gnd(gnd), .A(_1015__bF_buf0), .Y(_61_), .vdd(vdd), .B(_1966__bF_buf0), .C(_1974_), );
  NOR2X1 NOR2X1_116 (.gnd(gnd), .A(regs_10__8_), .Y(_1975_), .vdd(vdd), .B(_1966__bF_buf7), );
  AOI21X1 AOI21X1_105 (.gnd(gnd), .A(_1017__bF_buf0), .Y(_62_), .vdd(vdd), .B(_1966__bF_buf6), .C(_1975_), );
  NOR2X1 NOR2X1_117 (.gnd(gnd), .A(regs_10__9_), .Y(_1976_), .vdd(vdd), .B(_1966__bF_buf5), );
  AOI21X1 AOI21X1_106 (.gnd(gnd), .A(_1019__bF_buf0), .Y(_63_), .vdd(vdd), .B(_1966__bF_buf4), .C(_1976_), );
  NOR2X1 NOR2X1_118 (.gnd(gnd), .A(regs_10__10_), .Y(_1977_), .vdd(vdd), .B(_1966__bF_buf3), );
  AOI21X1 AOI21X1_107 (.gnd(gnd), .A(_1021__bF_buf0), .Y(_33_), .vdd(vdd), .B(_1966__bF_buf2), .C(_1977_), );
  NOR2X1 NOR2X1_119 (.gnd(gnd), .A(regs_10__11_), .Y(_1978_), .vdd(vdd), .B(_1966__bF_buf1), );
  AOI21X1 AOI21X1_108 (.gnd(gnd), .A(_1023__bF_buf0), .Y(_34_), .vdd(vdd), .B(_1966__bF_buf0), .C(_1978_), );
  NOR2X1 NOR2X1_120 (.gnd(gnd), .A(regs_10__12_), .Y(_1979_), .vdd(vdd), .B(_1966__bF_buf7), );
  AOI21X1 AOI21X1_109 (.gnd(gnd), .A(_1025__bF_buf0), .Y(_35_), .vdd(vdd), .B(_1966__bF_buf6), .C(_1979_), );
  NOR2X1 NOR2X1_121 (.gnd(gnd), .A(regs_10__13_), .Y(_1980_), .vdd(vdd), .B(_1966__bF_buf5), );
  AOI21X1 AOI21X1_110 (.gnd(gnd), .A(_1027__bF_buf0), .Y(_36_), .vdd(vdd), .B(_1966__bF_buf4), .C(_1980_), );
  NOR2X1 NOR2X1_122 (.gnd(gnd), .A(regs_10__14_), .Y(_1981_), .vdd(vdd), .B(_1966__bF_buf3), );
  AOI21X1 AOI21X1_111 (.gnd(gnd), .A(_1029__bF_buf0), .Y(_37_), .vdd(vdd), .B(_1966__bF_buf2), .C(_1981_), );
  NOR2X1 NOR2X1_123 (.gnd(gnd), .A(regs_10__15_), .Y(_1982_), .vdd(vdd), .B(_1966__bF_buf1), );
  AOI21X1 AOI21X1_112 (.gnd(gnd), .A(_1031__bF_buf0), .Y(_38_), .vdd(vdd), .B(_1966__bF_buf0), .C(_1982_), );
  NOR2X1 NOR2X1_124 (.gnd(gnd), .A(regs_10__16_), .Y(_1983_), .vdd(vdd), .B(_1966__bF_buf7), );
  AOI21X1 AOI21X1_113 (.gnd(gnd), .A(_1033__bF_buf0), .Y(_39_), .vdd(vdd), .B(_1966__bF_buf6), .C(_1983_), );
  NOR2X1 NOR2X1_125 (.gnd(gnd), .A(regs_10__17_), .Y(_1984_), .vdd(vdd), .B(_1966__bF_buf5), );
  AOI21X1 AOI21X1_114 (.gnd(gnd), .A(_1035__bF_buf0), .Y(_40_), .vdd(vdd), .B(_1966__bF_buf4), .C(_1984_), );
  NOR2X1 NOR2X1_126 (.gnd(gnd), .A(regs_10__18_), .Y(_1985_), .vdd(vdd), .B(_1966__bF_buf3), );
  AOI21X1 AOI21X1_115 (.gnd(gnd), .A(_1037__bF_buf0), .Y(_41_), .vdd(vdd), .B(_1966__bF_buf2), .C(_1985_), );
  NOR2X1 NOR2X1_127 (.gnd(gnd), .A(regs_10__19_), .Y(_1986_), .vdd(vdd), .B(_1966__bF_buf1), );
  AOI21X1 AOI21X1_116 (.gnd(gnd), .A(_1039__bF_buf0), .Y(_42_), .vdd(vdd), .B(_1966__bF_buf0), .C(_1986_), );
  NOR2X1 NOR2X1_128 (.gnd(gnd), .A(regs_10__20_), .Y(_1987_), .vdd(vdd), .B(_1966__bF_buf7), );
  AOI21X1 AOI21X1_117 (.gnd(gnd), .A(_1041__bF_buf0), .Y(_44_), .vdd(vdd), .B(_1966__bF_buf6), .C(_1987_), );
  NOR2X1 NOR2X1_129 (.gnd(gnd), .A(regs_10__21_), .Y(_1988_), .vdd(vdd), .B(_1966__bF_buf5), );
  AOI21X1 AOI21X1_118 (.gnd(gnd), .A(_1043__bF_buf0), .Y(_45_), .vdd(vdd), .B(_1966__bF_buf4), .C(_1988_), );
  NOR2X1 NOR2X1_130 (.gnd(gnd), .A(regs_10__22_), .Y(_1989_), .vdd(vdd), .B(_1966__bF_buf3), );
  AOI21X1 AOI21X1_119 (.gnd(gnd), .A(_1045__bF_buf0), .Y(_46_), .vdd(vdd), .B(_1966__bF_buf2), .C(_1989_), );
  NOR2X1 NOR2X1_131 (.gnd(gnd), .A(regs_10__23_), .Y(_1990_), .vdd(vdd), .B(_1966__bF_buf1), );
  AOI21X1 AOI21X1_120 (.gnd(gnd), .A(_1047__bF_buf0), .Y(_47_), .vdd(vdd), .B(_1966__bF_buf0), .C(_1990_), );
  NOR2X1 NOR2X1_132 (.gnd(gnd), .A(regs_10__24_), .Y(_1991_), .vdd(vdd), .B(_1966__bF_buf7), );
  AOI21X1 AOI21X1_121 (.gnd(gnd), .A(_1049__bF_buf0), .Y(_48_), .vdd(vdd), .B(_1966__bF_buf6), .C(_1991_), );
  NOR2X1 NOR2X1_133 (.gnd(gnd), .A(regs_10__25_), .Y(_1992_), .vdd(vdd), .B(_1966__bF_buf5), );
  AOI21X1 AOI21X1_122 (.gnd(gnd), .A(_1051__bF_buf0), .Y(_49_), .vdd(vdd), .B(_1966__bF_buf4), .C(_1992_), );
  NOR2X1 NOR2X1_134 (.gnd(gnd), .A(regs_10__26_), .Y(_1993_), .vdd(vdd), .B(_1966__bF_buf3), );
  AOI21X1 AOI21X1_123 (.gnd(gnd), .A(_1053__bF_buf0), .Y(_50_), .vdd(vdd), .B(_1966__bF_buf2), .C(_1993_), );
  NOR2X1 NOR2X1_135 (.gnd(gnd), .A(regs_10__27_), .Y(_1994_), .vdd(vdd), .B(_1966__bF_buf1), );
  AOI21X1 AOI21X1_124 (.gnd(gnd), .A(_1055__bF_buf0), .Y(_51_), .vdd(vdd), .B(_1966__bF_buf0), .C(_1994_), );
  NOR2X1 NOR2X1_136 (.gnd(gnd), .A(regs_10__28_), .Y(_1995_), .vdd(vdd), .B(_1966__bF_buf7), );
  AOI21X1 AOI21X1_125 (.gnd(gnd), .A(_1057__bF_buf0), .Y(_52_), .vdd(vdd), .B(_1966__bF_buf6), .C(_1995_), );
  NOR2X1 NOR2X1_137 (.gnd(gnd), .A(regs_10__29_), .Y(_1996_), .vdd(vdd), .B(_1966__bF_buf5), );
  AOI21X1 AOI21X1_126 (.gnd(gnd), .A(_1059__bF_buf0), .Y(_53_), .vdd(vdd), .B(_1966__bF_buf4), .C(_1996_), );
  NOR2X1 NOR2X1_138 (.gnd(gnd), .A(regs_10__30_), .Y(_1997_), .vdd(vdd), .B(_1966__bF_buf3), );
  AOI21X1 AOI21X1_127 (.gnd(gnd), .A(_1061__bF_buf0), .Y(_55_), .vdd(vdd), .B(_1966__bF_buf2), .C(_1997_), );
  NOR2X1 NOR2X1_139 (.gnd(gnd), .A(regs_10__31_), .Y(_1998_), .vdd(vdd), .B(_1966__bF_buf1), );
  AOI21X1 AOI21X1_128 (.gnd(gnd), .A(_1063__bF_buf0), .Y(_56_), .vdd(vdd), .B(_1966__bF_buf0), .C(_1998_), );
  INVX2 INVX2_225 (.gnd(gnd), .A(regs_9__0_), .Y(_1999_), .vdd(vdd), );
  NOR2X1 NOR2X1_140 (.gnd(gnd), .A(_1901__bF_buf3), .Y(_2000_), .vdd(vdd), .B(_1070__bF_buf7), );
  NAND2X1 NAND2X1_227 (.gnd(gnd), .A(wdata[0]), .Y(_2001_), .vdd(vdd), .B(_2000__bF_buf7), );
  OAI21X1 OAI21X1_473 (.gnd(gnd), .A(_1999_), .Y(_960_), .vdd(vdd), .B(_2000__bF_buf6), .C(_2001_), );
  INVX2 INVX2_226 (.gnd(gnd), .A(regs_9__1_), .Y(_2002_), .vdd(vdd), );
  NAND2X1 NAND2X1_228 (.gnd(gnd), .A(wdata[1]), .Y(_2003_), .vdd(vdd), .B(_2000__bF_buf5), );
  OAI21X1 OAI21X1_474 (.gnd(gnd), .A(_2002_), .Y(_971_), .vdd(vdd), .B(_2000__bF_buf4), .C(_2003_), );
  INVX2 INVX2_227 (.gnd(gnd), .A(regs_9__2_), .Y(_2004_), .vdd(vdd), );
  NAND2X1 NAND2X1_229 (.gnd(gnd), .A(wdata[2]), .Y(_2005_), .vdd(vdd), .B(_2000__bF_buf3), );
  OAI21X1 OAI21X1_475 (.gnd(gnd), .A(_2004_), .Y(_982_), .vdd(vdd), .B(_2000__bF_buf2), .C(_2005_), );
  INVX2 INVX2_228 (.gnd(gnd), .A(regs_9__3_), .Y(_2006_), .vdd(vdd), );
  NAND2X1 NAND2X1_230 (.gnd(gnd), .A(wdata[3]), .Y(_2007_), .vdd(vdd), .B(_2000__bF_buf1), );
  OAI21X1 OAI21X1_476 (.gnd(gnd), .A(_2006_), .Y(_985_), .vdd(vdd), .B(_2000__bF_buf0), .C(_2007_), );
  INVX2 INVX2_229 (.gnd(gnd), .A(regs_9__4_), .Y(_2008_), .vdd(vdd), );
  NAND2X1 NAND2X1_231 (.gnd(gnd), .A(wdata[4]), .Y(_2009_), .vdd(vdd), .B(_2000__bF_buf7), );
  OAI21X1 OAI21X1_477 (.gnd(gnd), .A(_2008_), .Y(_986_), .vdd(vdd), .B(_2000__bF_buf6), .C(_2009_), );
  INVX2 INVX2_230 (.gnd(gnd), .A(regs_9__5_), .Y(_2010_), .vdd(vdd), );
  NAND2X1 NAND2X1_232 (.gnd(gnd), .A(wdata[5]), .Y(_2011_), .vdd(vdd), .B(_2000__bF_buf5), );
  OAI21X1 OAI21X1_478 (.gnd(gnd), .A(_2010_), .Y(_987_), .vdd(vdd), .B(_2000__bF_buf4), .C(_2011_), );
  INVX2 INVX2_231 (.gnd(gnd), .A(regs_9__6_), .Y(_2012_), .vdd(vdd), );
  NAND2X1 NAND2X1_233 (.gnd(gnd), .A(wdata[6]), .Y(_2013_), .vdd(vdd), .B(_2000__bF_buf3), );
  OAI21X1 OAI21X1_479 (.gnd(gnd), .A(_2012_), .Y(_988_), .vdd(vdd), .B(_2000__bF_buf2), .C(_2013_), );
  INVX2 INVX2_232 (.gnd(gnd), .A(regs_9__7_), .Y(_2014_), .vdd(vdd), );
  NAND2X1 NAND2X1_234 (.gnd(gnd), .A(wdata[7]), .Y(_2015_), .vdd(vdd), .B(_2000__bF_buf1), );
  OAI21X1 OAI21X1_480 (.gnd(gnd), .A(_2014_), .Y(_989_), .vdd(vdd), .B(_2000__bF_buf0), .C(_2015_), );
  INVX2 INVX2_233 (.gnd(gnd), .A(regs_9__8_), .Y(_2016_), .vdd(vdd), );
  NAND2X1 NAND2X1_235 (.gnd(gnd), .A(wdata[8]), .Y(_2017_), .vdd(vdd), .B(_2000__bF_buf7), );
  OAI21X1 OAI21X1_481 (.gnd(gnd), .A(_2016_), .Y(_990_), .vdd(vdd), .B(_2000__bF_buf6), .C(_2017_), );
  INVX2 INVX2_234 (.gnd(gnd), .A(regs_9__9_), .Y(_2018_), .vdd(vdd), );
  NAND2X1 NAND2X1_236 (.gnd(gnd), .A(wdata[9]), .Y(_2019_), .vdd(vdd), .B(_2000__bF_buf5), );
  OAI21X1 OAI21X1_482 (.gnd(gnd), .A(_2018_), .Y(_991_), .vdd(vdd), .B(_2000__bF_buf4), .C(_2019_), );
  INVX2 INVX2_235 (.gnd(gnd), .A(regs_9__10_), .Y(_2020_), .vdd(vdd), );
  NAND2X1 NAND2X1_237 (.gnd(gnd), .A(wdata[10]), .Y(_2021_), .vdd(vdd), .B(_2000__bF_buf3), );
  OAI21X1 OAI21X1_483 (.gnd(gnd), .A(_2020_), .Y(_961_), .vdd(vdd), .B(_2000__bF_buf2), .C(_2021_), );
  INVX2 INVX2_236 (.gnd(gnd), .A(regs_9__11_), .Y(_2022_), .vdd(vdd), );
  NAND2X1 NAND2X1_238 (.gnd(gnd), .A(wdata[11]), .Y(_2023_), .vdd(vdd), .B(_2000__bF_buf1), );
  OAI21X1 OAI21X1_484 (.gnd(gnd), .A(_2022_), .Y(_962_), .vdd(vdd), .B(_2000__bF_buf0), .C(_2023_), );
  INVX2 INVX2_237 (.gnd(gnd), .A(regs_9__12_), .Y(_2024_), .vdd(vdd), );
  NAND2X1 NAND2X1_239 (.gnd(gnd), .A(wdata[12]), .Y(_2025_), .vdd(vdd), .B(_2000__bF_buf7), );
  OAI21X1 OAI21X1_485 (.gnd(gnd), .A(_2024_), .Y(_963_), .vdd(vdd), .B(_2000__bF_buf6), .C(_2025_), );
  INVX2 INVX2_238 (.gnd(gnd), .A(regs_9__13_), .Y(_2026_), .vdd(vdd), );
  NAND2X1 NAND2X1_240 (.gnd(gnd), .A(wdata[13]), .Y(_2027_), .vdd(vdd), .B(_2000__bF_buf5), );
  OAI21X1 OAI21X1_486 (.gnd(gnd), .A(_2026_), .Y(_964_), .vdd(vdd), .B(_2000__bF_buf4), .C(_2027_), );
  INVX2 INVX2_239 (.gnd(gnd), .A(regs_9__14_), .Y(_2028_), .vdd(vdd), );
  NAND2X1 NAND2X1_241 (.gnd(gnd), .A(wdata[14]), .Y(_2029_), .vdd(vdd), .B(_2000__bF_buf3), );
  OAI21X1 OAI21X1_487 (.gnd(gnd), .A(_2028_), .Y(_965_), .vdd(vdd), .B(_2000__bF_buf2), .C(_2029_), );
  INVX2 INVX2_240 (.gnd(gnd), .A(regs_9__15_), .Y(_2030_), .vdd(vdd), );
  NAND2X1 NAND2X1_242 (.gnd(gnd), .A(wdata[15]), .Y(_2031_), .vdd(vdd), .B(_2000__bF_buf1), );
  OAI21X1 OAI21X1_488 (.gnd(gnd), .A(_2030_), .Y(_966_), .vdd(vdd), .B(_2000__bF_buf0), .C(_2031_), );
  INVX2 INVX2_241 (.gnd(gnd), .A(regs_9__16_), .Y(_2032_), .vdd(vdd), );
  NAND2X1 NAND2X1_243 (.gnd(gnd), .A(wdata[16]), .Y(_2033_), .vdd(vdd), .B(_2000__bF_buf7), );
  OAI21X1 OAI21X1_489 (.gnd(gnd), .A(_2032_), .Y(_967_), .vdd(vdd), .B(_2000__bF_buf6), .C(_2033_), );
  INVX2 INVX2_242 (.gnd(gnd), .A(regs_9__17_), .Y(_2034_), .vdd(vdd), );
  NAND2X1 NAND2X1_244 (.gnd(gnd), .A(wdata[17]), .Y(_2035_), .vdd(vdd), .B(_2000__bF_buf5), );
  OAI21X1 OAI21X1_490 (.gnd(gnd), .A(_2034_), .Y(_968_), .vdd(vdd), .B(_2000__bF_buf4), .C(_2035_), );
  INVX2 INVX2_243 (.gnd(gnd), .A(regs_9__18_), .Y(_2036_), .vdd(vdd), );
  NAND2X1 NAND2X1_245 (.gnd(gnd), .A(wdata[18]), .Y(_2037_), .vdd(vdd), .B(_2000__bF_buf3), );
  OAI21X1 OAI21X1_491 (.gnd(gnd), .A(_2036_), .Y(_969_), .vdd(vdd), .B(_2000__bF_buf2), .C(_2037_), );
  INVX2 INVX2_244 (.gnd(gnd), .A(regs_9__19_), .Y(_2038_), .vdd(vdd), );
  NAND2X1 NAND2X1_246 (.gnd(gnd), .A(wdata[19]), .Y(_2039_), .vdd(vdd), .B(_2000__bF_buf1), );
  OAI21X1 OAI21X1_492 (.gnd(gnd), .A(_2038_), .Y(_970_), .vdd(vdd), .B(_2000__bF_buf0), .C(_2039_), );
  INVX2 INVX2_245 (.gnd(gnd), .A(regs_9__20_), .Y(_2040_), .vdd(vdd), );
  NAND2X1 NAND2X1_247 (.gnd(gnd), .A(wdata[20]), .Y(_2041_), .vdd(vdd), .B(_2000__bF_buf7), );
  OAI21X1 OAI21X1_493 (.gnd(gnd), .A(_2040_), .Y(_972_), .vdd(vdd), .B(_2000__bF_buf6), .C(_2041_), );
  INVX2 INVX2_246 (.gnd(gnd), .A(regs_9__21_), .Y(_2042_), .vdd(vdd), );
  NAND2X1 NAND2X1_248 (.gnd(gnd), .A(wdata[21]), .Y(_2043_), .vdd(vdd), .B(_2000__bF_buf5), );
  OAI21X1 OAI21X1_494 (.gnd(gnd), .A(_2042_), .Y(_973_), .vdd(vdd), .B(_2000__bF_buf4), .C(_2043_), );
  INVX2 INVX2_247 (.gnd(gnd), .A(regs_9__22_), .Y(_2044_), .vdd(vdd), );
  NAND2X1 NAND2X1_249 (.gnd(gnd), .A(wdata[22]), .Y(_2045_), .vdd(vdd), .B(_2000__bF_buf3), );
  OAI21X1 OAI21X1_495 (.gnd(gnd), .A(_2044_), .Y(_974_), .vdd(vdd), .B(_2000__bF_buf2), .C(_2045_), );
  INVX2 INVX2_248 (.gnd(gnd), .A(regs_9__23_), .Y(_2046_), .vdd(vdd), );
  NAND2X1 NAND2X1_250 (.gnd(gnd), .A(wdata[23]), .Y(_2047_), .vdd(vdd), .B(_2000__bF_buf1), );
  OAI21X1 OAI21X1_496 (.gnd(gnd), .A(_2046_), .Y(_975_), .vdd(vdd), .B(_2000__bF_buf0), .C(_2047_), );
  INVX2 INVX2_249 (.gnd(gnd), .A(regs_9__24_), .Y(_2048_), .vdd(vdd), );
  NAND2X1 NAND2X1_251 (.gnd(gnd), .A(wdata[24]), .Y(_2049_), .vdd(vdd), .B(_2000__bF_buf7), );
  OAI21X1 OAI21X1_497 (.gnd(gnd), .A(_2048_), .Y(_976_), .vdd(vdd), .B(_2000__bF_buf6), .C(_2049_), );
  INVX2 INVX2_250 (.gnd(gnd), .A(regs_9__25_), .Y(_2050_), .vdd(vdd), );
  NAND2X1 NAND2X1_252 (.gnd(gnd), .A(wdata[25]), .Y(_2051_), .vdd(vdd), .B(_2000__bF_buf5), );
  OAI21X1 OAI21X1_498 (.gnd(gnd), .A(_2050_), .Y(_977_), .vdd(vdd), .B(_2000__bF_buf4), .C(_2051_), );
  INVX2 INVX2_251 (.gnd(gnd), .A(regs_9__26_), .Y(_2052_), .vdd(vdd), );
  NAND2X1 NAND2X1_253 (.gnd(gnd), .A(wdata[26]), .Y(_2053_), .vdd(vdd), .B(_2000__bF_buf3), );
  OAI21X1 OAI21X1_499 (.gnd(gnd), .A(_2052_), .Y(_978_), .vdd(vdd), .B(_2000__bF_buf2), .C(_2053_), );
  INVX2 INVX2_252 (.gnd(gnd), .A(regs_9__27_), .Y(_2054_), .vdd(vdd), );
  NAND2X1 NAND2X1_254 (.gnd(gnd), .A(wdata[27]), .Y(_2055_), .vdd(vdd), .B(_2000__bF_buf1), );
  OAI21X1 OAI21X1_500 (.gnd(gnd), .A(_2054_), .Y(_979_), .vdd(vdd), .B(_2000__bF_buf0), .C(_2055_), );
  INVX2 INVX2_253 (.gnd(gnd), .A(regs_9__28_), .Y(_2056_), .vdd(vdd), );
  NAND2X1 NAND2X1_255 (.gnd(gnd), .A(wdata[28]), .Y(_2057_), .vdd(vdd), .B(_2000__bF_buf7), );
  OAI21X1 OAI21X1_501 (.gnd(gnd), .A(_2056_), .Y(_980_), .vdd(vdd), .B(_2000__bF_buf6), .C(_2057_), );
  INVX2 INVX2_254 (.gnd(gnd), .A(regs_9__29_), .Y(_2058_), .vdd(vdd), );
  NAND2X1 NAND2X1_256 (.gnd(gnd), .A(wdata[29]), .Y(_2059_), .vdd(vdd), .B(_2000__bF_buf5), );
  OAI21X1 OAI21X1_502 (.gnd(gnd), .A(_2058_), .Y(_981_), .vdd(vdd), .B(_2000__bF_buf4), .C(_2059_), );
  INVX2 INVX2_255 (.gnd(gnd), .A(regs_9__30_), .Y(_2060_), .vdd(vdd), );
  NAND2X1 NAND2X1_257 (.gnd(gnd), .A(wdata[30]), .Y(_2061_), .vdd(vdd), .B(_2000__bF_buf3), );
  OAI21X1 OAI21X1_503 (.gnd(gnd), .A(_2060_), .Y(_983_), .vdd(vdd), .B(_2000__bF_buf2), .C(_2061_), );
  INVX2 INVX2_256 (.gnd(gnd), .A(regs_9__31_), .Y(_2062_), .vdd(vdd), );
  NAND2X1 NAND2X1_258 (.gnd(gnd), .A(wdata[31]), .Y(_2063_), .vdd(vdd), .B(_2000__bF_buf1), );
  OAI21X1 OAI21X1_504 (.gnd(gnd), .A(_2062_), .Y(_984_), .vdd(vdd), .B(_2000__bF_buf0), .C(_2063_), );
  OR2X2 OR2X2_8 (.gnd(gnd), .A(_1901__bF_buf2), .Y(_2064_), .vdd(vdd), .B(_1104__bF_buf7), );
  OAI21X1 OAI21X1_505 (.gnd(gnd), .A(_1901__bF_buf1), .Y(_2065_), .vdd(vdd), .B(_1104__bF_buf6), .C(regs_8__0_), );
  OAI21X1 OAI21X1_506 (.gnd(gnd), .A(_2064__bF_buf4), .Y(_928_), .vdd(vdd), .B(_992__bF_buf0), .C(_2065_), );
  OAI21X1 OAI21X1_507 (.gnd(gnd), .A(_1901__bF_buf0), .Y(_2066_), .vdd(vdd), .B(_1104__bF_buf5), .C(regs_8__1_), );
  OAI21X1 OAI21X1_508 (.gnd(gnd), .A(_2064__bF_buf3), .Y(_939_), .vdd(vdd), .B(_1003__bF_buf0), .C(_2066_), );
  OAI21X1 OAI21X1_509 (.gnd(gnd), .A(_1901__bF_buf5), .Y(_2067_), .vdd(vdd), .B(_1104__bF_buf4), .C(regs_8__2_), );
  OAI21X1 OAI21X1_510 (.gnd(gnd), .A(_2064__bF_buf2), .Y(_950_), .vdd(vdd), .B(_1005__bF_buf0), .C(_2067_), );
  OAI21X1 OAI21X1_511 (.gnd(gnd), .A(_1901__bF_buf4), .Y(_2068_), .vdd(vdd), .B(_1104__bF_buf3), .C(regs_8__3_), );
  OAI21X1 OAI21X1_512 (.gnd(gnd), .A(_2064__bF_buf1), .Y(_953_), .vdd(vdd), .B(_1007__bF_buf0), .C(_2068_), );
  OAI21X1 OAI21X1_513 (.gnd(gnd), .A(_1901__bF_buf3), .Y(_2069_), .vdd(vdd), .B(_1104__bF_buf2), .C(regs_8__4_), );
  OAI21X1 OAI21X1_514 (.gnd(gnd), .A(_2064__bF_buf0), .Y(_954_), .vdd(vdd), .B(_1009__bF_buf3), .C(_2069_), );
  OAI21X1 OAI21X1_515 (.gnd(gnd), .A(_1901__bF_buf2), .Y(_2070_), .vdd(vdd), .B(_1104__bF_buf1), .C(regs_8__5_), );
  OAI21X1 OAI21X1_516 (.gnd(gnd), .A(_2064__bF_buf4), .Y(_955_), .vdd(vdd), .B(_1011__bF_buf3), .C(_2070_), );
  OAI21X1 OAI21X1_517 (.gnd(gnd), .A(_1901__bF_buf1), .Y(_2071_), .vdd(vdd), .B(_1104__bF_buf0), .C(regs_8__6_), );
  OAI21X1 OAI21X1_518 (.gnd(gnd), .A(_2064__bF_buf3), .Y(_956_), .vdd(vdd), .B(_1013__bF_buf3), .C(_2071_), );
  OAI21X1 OAI21X1_519 (.gnd(gnd), .A(_1901__bF_buf0), .Y(_2072_), .vdd(vdd), .B(_1104__bF_buf14), .C(regs_8__7_), );
  OAI21X1 OAI21X1_520 (.gnd(gnd), .A(_2064__bF_buf2), .Y(_957_), .vdd(vdd), .B(_1015__bF_buf3), .C(_2072_), );
  OAI21X1 OAI21X1_521 (.gnd(gnd), .A(_1901__bF_buf5), .Y(_2073_), .vdd(vdd), .B(_1104__bF_buf13), .C(regs_8__8_), );
  OAI21X1 OAI21X1_522 (.gnd(gnd), .A(_2064__bF_buf1), .Y(_958_), .vdd(vdd), .B(_1017__bF_buf3), .C(_2073_), );
  OAI21X1 OAI21X1_523 (.gnd(gnd), .A(_1901__bF_buf4), .Y(_2074_), .vdd(vdd), .B(_1104__bF_buf12), .C(regs_8__9_), );
  OAI21X1 OAI21X1_524 (.gnd(gnd), .A(_2064__bF_buf0), .Y(_959_), .vdd(vdd), .B(_1019__bF_buf3), .C(_2074_), );
  OAI21X1 OAI21X1_525 (.gnd(gnd), .A(_1901__bF_buf3), .Y(_2075_), .vdd(vdd), .B(_1104__bF_buf11), .C(regs_8__10_), );
  OAI21X1 OAI21X1_526 (.gnd(gnd), .A(_2064__bF_buf4), .Y(_929_), .vdd(vdd), .B(_1021__bF_buf3), .C(_2075_), );
  OAI21X1 OAI21X1_527 (.gnd(gnd), .A(_1901__bF_buf2), .Y(_2076_), .vdd(vdd), .B(_1104__bF_buf10), .C(regs_8__11_), );
  OAI21X1 OAI21X1_528 (.gnd(gnd), .A(_2064__bF_buf3), .Y(_930_), .vdd(vdd), .B(_1023__bF_buf3), .C(_2076_), );
  OAI21X1 OAI21X1_529 (.gnd(gnd), .A(_1901__bF_buf1), .Y(_2077_), .vdd(vdd), .B(_1104__bF_buf9), .C(regs_8__12_), );
  OAI21X1 OAI21X1_530 (.gnd(gnd), .A(_2064__bF_buf2), .Y(_931_), .vdd(vdd), .B(_1025__bF_buf3), .C(_2077_), );
  OAI21X1 OAI21X1_531 (.gnd(gnd), .A(_1901__bF_buf0), .Y(_2078_), .vdd(vdd), .B(_1104__bF_buf8), .C(regs_8__13_), );
  OAI21X1 OAI21X1_532 (.gnd(gnd), .A(_2064__bF_buf1), .Y(_932_), .vdd(vdd), .B(_1027__bF_buf3), .C(_2078_), );
  OAI21X1 OAI21X1_533 (.gnd(gnd), .A(_1901__bF_buf5), .Y(_2079_), .vdd(vdd), .B(_1104__bF_buf7), .C(regs_8__14_), );
  OAI21X1 OAI21X1_534 (.gnd(gnd), .A(_2064__bF_buf0), .Y(_933_), .vdd(vdd), .B(_1029__bF_buf3), .C(_2079_), );
  OAI21X1 OAI21X1_535 (.gnd(gnd), .A(_1901__bF_buf4), .Y(_2080_), .vdd(vdd), .B(_1104__bF_buf6), .C(regs_8__15_), );
  OAI21X1 OAI21X1_536 (.gnd(gnd), .A(_2064__bF_buf4), .Y(_934_), .vdd(vdd), .B(_1031__bF_buf3), .C(_2080_), );
  OAI21X1 OAI21X1_537 (.gnd(gnd), .A(_1901__bF_buf3), .Y(_2081_), .vdd(vdd), .B(_1104__bF_buf5), .C(regs_8__16_), );
  OAI21X1 OAI21X1_538 (.gnd(gnd), .A(_2064__bF_buf3), .Y(_935_), .vdd(vdd), .B(_1033__bF_buf3), .C(_2081_), );
  OAI21X1 OAI21X1_539 (.gnd(gnd), .A(_1901__bF_buf2), .Y(_2082_), .vdd(vdd), .B(_1104__bF_buf4), .C(regs_8__17_), );
  OAI21X1 OAI21X1_540 (.gnd(gnd), .A(_2064__bF_buf2), .Y(_936_), .vdd(vdd), .B(_1035__bF_buf3), .C(_2082_), );
  OAI21X1 OAI21X1_541 (.gnd(gnd), .A(_1901__bF_buf1), .Y(_2083_), .vdd(vdd), .B(_1104__bF_buf3), .C(regs_8__18_), );
  OAI21X1 OAI21X1_542 (.gnd(gnd), .A(_2064__bF_buf1), .Y(_937_), .vdd(vdd), .B(_1037__bF_buf3), .C(_2083_), );
  OAI21X1 OAI21X1_543 (.gnd(gnd), .A(_1901__bF_buf0), .Y(_2084_), .vdd(vdd), .B(_1104__bF_buf2), .C(regs_8__19_), );
  OAI21X1 OAI21X1_544 (.gnd(gnd), .A(_2064__bF_buf0), .Y(_938_), .vdd(vdd), .B(_1039__bF_buf3), .C(_2084_), );
  OAI21X1 OAI21X1_545 (.gnd(gnd), .A(_1901__bF_buf5), .Y(_2085_), .vdd(vdd), .B(_1104__bF_buf1), .C(regs_8__20_), );
  OAI21X1 OAI21X1_546 (.gnd(gnd), .A(_2064__bF_buf4), .Y(_940_), .vdd(vdd), .B(_1041__bF_buf3), .C(_2085_), );
  OAI21X1 OAI21X1_547 (.gnd(gnd), .A(_1901__bF_buf4), .Y(_2086_), .vdd(vdd), .B(_1104__bF_buf0), .C(regs_8__21_), );
  OAI21X1 OAI21X1_548 (.gnd(gnd), .A(_2064__bF_buf3), .Y(_941_), .vdd(vdd), .B(_1043__bF_buf3), .C(_2086_), );
  OAI21X1 OAI21X1_549 (.gnd(gnd), .A(_1901__bF_buf3), .Y(_2087_), .vdd(vdd), .B(_1104__bF_buf14), .C(regs_8__22_), );
  OAI21X1 OAI21X1_550 (.gnd(gnd), .A(_2064__bF_buf2), .Y(_942_), .vdd(vdd), .B(_1045__bF_buf3), .C(_2087_), );
  OAI21X1 OAI21X1_551 (.gnd(gnd), .A(_1901__bF_buf2), .Y(_2088_), .vdd(vdd), .B(_1104__bF_buf13), .C(regs_8__23_), );
  OAI21X1 OAI21X1_552 (.gnd(gnd), .A(_2064__bF_buf1), .Y(_943_), .vdd(vdd), .B(_1047__bF_buf3), .C(_2088_), );
  OAI21X1 OAI21X1_553 (.gnd(gnd), .A(_1901__bF_buf1), .Y(_2089_), .vdd(vdd), .B(_1104__bF_buf12), .C(regs_8__24_), );
  OAI21X1 OAI21X1_554 (.gnd(gnd), .A(_2064__bF_buf0), .Y(_944_), .vdd(vdd), .B(_1049__bF_buf3), .C(_2089_), );
  OAI21X1 OAI21X1_555 (.gnd(gnd), .A(_1901__bF_buf0), .Y(_2090_), .vdd(vdd), .B(_1104__bF_buf11), .C(regs_8__25_), );
  OAI21X1 OAI21X1_556 (.gnd(gnd), .A(_2064__bF_buf4), .Y(_945_), .vdd(vdd), .B(_1051__bF_buf3), .C(_2090_), );
  OAI21X1 OAI21X1_557 (.gnd(gnd), .A(_1901__bF_buf5), .Y(_2091_), .vdd(vdd), .B(_1104__bF_buf10), .C(regs_8__26_), );
  OAI21X1 OAI21X1_558 (.gnd(gnd), .A(_2064__bF_buf3), .Y(_946_), .vdd(vdd), .B(_1053__bF_buf3), .C(_2091_), );
  OAI21X1 OAI21X1_559 (.gnd(gnd), .A(_1901__bF_buf4), .Y(_2092_), .vdd(vdd), .B(_1104__bF_buf9), .C(regs_8__27_), );
  OAI21X1 OAI21X1_560 (.gnd(gnd), .A(_2064__bF_buf2), .Y(_947_), .vdd(vdd), .B(_1055__bF_buf3), .C(_2092_), );
  OAI21X1 OAI21X1_561 (.gnd(gnd), .A(_1901__bF_buf3), .Y(_2093_), .vdd(vdd), .B(_1104__bF_buf8), .C(regs_8__28_), );
  OAI21X1 OAI21X1_562 (.gnd(gnd), .A(_2064__bF_buf1), .Y(_948_), .vdd(vdd), .B(_1057__bF_buf3), .C(_2093_), );
  OAI21X1 OAI21X1_563 (.gnd(gnd), .A(_1901__bF_buf2), .Y(_2094_), .vdd(vdd), .B(_1104__bF_buf7), .C(regs_8__29_), );
  OAI21X1 OAI21X1_564 (.gnd(gnd), .A(_2064__bF_buf0), .Y(_949_), .vdd(vdd), .B(_1059__bF_buf3), .C(_2094_), );
  OAI21X1 OAI21X1_565 (.gnd(gnd), .A(_1901__bF_buf1), .Y(_2095_), .vdd(vdd), .B(_1104__bF_buf6), .C(regs_8__30_), );
  OAI21X1 OAI21X1_566 (.gnd(gnd), .A(_2064__bF_buf4), .Y(_951_), .vdd(vdd), .B(_1061__bF_buf3), .C(_2095_), );
  OAI21X1 OAI21X1_567 (.gnd(gnd), .A(_1901__bF_buf0), .Y(_2096_), .vdd(vdd), .B(_1104__bF_buf5), .C(regs_8__31_), );
  OAI21X1 OAI21X1_568 (.gnd(gnd), .A(_2064__bF_buf3), .Y(_952_), .vdd(vdd), .B(_1063__bF_buf3), .C(_2096_), );
  INVX2 INVX2_257 (.gnd(gnd), .A(regs_7__0_), .Y(_2097_), .vdd(vdd), );
  NAND2X1 NAND2X1_259 (.gnd(gnd), .A(waddr[4]), .Y(_2098_), .vdd(vdd), .B(waddr[3]), );
  NOR2X1 NOR2X1_141 (.gnd(gnd), .A(waddr[2]), .Y(_2099_), .vdd(vdd), .B(_2098_), );
  INVX8 INVX8_1 (.gnd(gnd), .A(_2099_), .Y(_2100_), .vdd(vdd), );
  NOR2X1 NOR2X1_142 (.gnd(gnd), .A(_1142__bF_buf1), .Y(_2101_), .vdd(vdd), .B(_2100__bF_buf8), );
  NAND2X1 NAND2X1_260 (.gnd(gnd), .A(wdata[0]), .Y(_2102_), .vdd(vdd), .B(_2101__bF_buf7), );
  OAI21X1 OAI21X1_569 (.gnd(gnd), .A(_2097_), .Y(_896_), .vdd(vdd), .B(_2101__bF_buf6), .C(_2102_), );
  INVX2 INVX2_258 (.gnd(gnd), .A(regs_7__1_), .Y(_2103_), .vdd(vdd), );
  NAND2X1 NAND2X1_261 (.gnd(gnd), .A(wdata[1]), .Y(_2104_), .vdd(vdd), .B(_2101__bF_buf5), );
  OAI21X1 OAI21X1_570 (.gnd(gnd), .A(_2103_), .Y(_907_), .vdd(vdd), .B(_2101__bF_buf4), .C(_2104_), );
  INVX2 INVX2_259 (.gnd(gnd), .A(regs_7__2_), .Y(_2105_), .vdd(vdd), );
  NAND2X1 NAND2X1_262 (.gnd(gnd), .A(wdata[2]), .Y(_2106_), .vdd(vdd), .B(_2101__bF_buf3), );
  OAI21X1 OAI21X1_571 (.gnd(gnd), .A(_2105_), .Y(_918_), .vdd(vdd), .B(_2101__bF_buf2), .C(_2106_), );
  INVX2 INVX2_260 (.gnd(gnd), .A(regs_7__3_), .Y(_2107_), .vdd(vdd), );
  NAND2X1 NAND2X1_263 (.gnd(gnd), .A(wdata[3]), .Y(_2108_), .vdd(vdd), .B(_2101__bF_buf1), );
  OAI21X1 OAI21X1_572 (.gnd(gnd), .A(_2107_), .Y(_921_), .vdd(vdd), .B(_2101__bF_buf0), .C(_2108_), );
  INVX2 INVX2_261 (.gnd(gnd), .A(regs_7__4_), .Y(_2109_), .vdd(vdd), );
  NAND2X1 NAND2X1_264 (.gnd(gnd), .A(wdata[4]), .Y(_2110_), .vdd(vdd), .B(_2101__bF_buf7), );
  OAI21X1 OAI21X1_573 (.gnd(gnd), .A(_2109_), .Y(_922_), .vdd(vdd), .B(_2101__bF_buf6), .C(_2110_), );
  INVX2 INVX2_262 (.gnd(gnd), .A(regs_7__5_), .Y(_2111_), .vdd(vdd), );
  NAND2X1 NAND2X1_265 (.gnd(gnd), .A(wdata[5]), .Y(_2112_), .vdd(vdd), .B(_2101__bF_buf5), );
  OAI21X1 OAI21X1_574 (.gnd(gnd), .A(_2111_), .Y(_923_), .vdd(vdd), .B(_2101__bF_buf4), .C(_2112_), );
  INVX2 INVX2_263 (.gnd(gnd), .A(regs_7__6_), .Y(_2113_), .vdd(vdd), );
  NAND2X1 NAND2X1_266 (.gnd(gnd), .A(wdata[6]), .Y(_2114_), .vdd(vdd), .B(_2101__bF_buf3), );
  OAI21X1 OAI21X1_575 (.gnd(gnd), .A(_2113_), .Y(_924_), .vdd(vdd), .B(_2101__bF_buf2), .C(_2114_), );
  INVX2 INVX2_264 (.gnd(gnd), .A(regs_7__7_), .Y(_2115_), .vdd(vdd), );
  NAND2X1 NAND2X1_267 (.gnd(gnd), .A(wdata[7]), .Y(_2116_), .vdd(vdd), .B(_2101__bF_buf1), );
  OAI21X1 OAI21X1_576 (.gnd(gnd), .A(_2115_), .Y(_925_), .vdd(vdd), .B(_2101__bF_buf0), .C(_2116_), );
  INVX2 INVX2_265 (.gnd(gnd), .A(regs_7__8_), .Y(_2117_), .vdd(vdd), );
  NAND2X1 NAND2X1_268 (.gnd(gnd), .A(wdata[8]), .Y(_2118_), .vdd(vdd), .B(_2101__bF_buf7), );
  OAI21X1 OAI21X1_577 (.gnd(gnd), .A(_2117_), .Y(_926_), .vdd(vdd), .B(_2101__bF_buf6), .C(_2118_), );
  INVX2 INVX2_266 (.gnd(gnd), .A(regs_7__9_), .Y(_2119_), .vdd(vdd), );
  NAND2X1 NAND2X1_269 (.gnd(gnd), .A(wdata[9]), .Y(_2120_), .vdd(vdd), .B(_2101__bF_buf5), );
  OAI21X1 OAI21X1_578 (.gnd(gnd), .A(_2119_), .Y(_927_), .vdd(vdd), .B(_2101__bF_buf4), .C(_2120_), );
  INVX2 INVX2_267 (.gnd(gnd), .A(regs_7__10_), .Y(_2121_), .vdd(vdd), );
  NAND2X1 NAND2X1_270 (.gnd(gnd), .A(wdata[10]), .Y(_2122_), .vdd(vdd), .B(_2101__bF_buf3), );
  OAI21X1 OAI21X1_579 (.gnd(gnd), .A(_2121_), .Y(_897_), .vdd(vdd), .B(_2101__bF_buf2), .C(_2122_), );
  INVX2 INVX2_268 (.gnd(gnd), .A(regs_7__11_), .Y(_2123_), .vdd(vdd), );
  NAND2X1 NAND2X1_271 (.gnd(gnd), .A(wdata[11]), .Y(_2124_), .vdd(vdd), .B(_2101__bF_buf1), );
  OAI21X1 OAI21X1_580 (.gnd(gnd), .A(_2123_), .Y(_898_), .vdd(vdd), .B(_2101__bF_buf0), .C(_2124_), );
  INVX2 INVX2_269 (.gnd(gnd), .A(regs_7__12_), .Y(_2125_), .vdd(vdd), );
  NAND2X1 NAND2X1_272 (.gnd(gnd), .A(wdata[12]), .Y(_2126_), .vdd(vdd), .B(_2101__bF_buf7), );
  OAI21X1 OAI21X1_581 (.gnd(gnd), .A(_2125_), .Y(_899_), .vdd(vdd), .B(_2101__bF_buf6), .C(_2126_), );
  INVX2 INVX2_270 (.gnd(gnd), .A(regs_7__13_), .Y(_2127_), .vdd(vdd), );
  NAND2X1 NAND2X1_273 (.gnd(gnd), .A(wdata[13]), .Y(_2128_), .vdd(vdd), .B(_2101__bF_buf5), );
  OAI21X1 OAI21X1_582 (.gnd(gnd), .A(_2127_), .Y(_900_), .vdd(vdd), .B(_2101__bF_buf4), .C(_2128_), );
  INVX2 INVX2_271 (.gnd(gnd), .A(regs_7__14_), .Y(_2129_), .vdd(vdd), );
  NAND2X1 NAND2X1_274 (.gnd(gnd), .A(wdata[14]), .Y(_2130_), .vdd(vdd), .B(_2101__bF_buf3), );
  OAI21X1 OAI21X1_583 (.gnd(gnd), .A(_2129_), .Y(_901_), .vdd(vdd), .B(_2101__bF_buf2), .C(_2130_), );
  INVX2 INVX2_272 (.gnd(gnd), .A(regs_7__15_), .Y(_2131_), .vdd(vdd), );
  NAND2X1 NAND2X1_275 (.gnd(gnd), .A(wdata[15]), .Y(_2132_), .vdd(vdd), .B(_2101__bF_buf1), );
  OAI21X1 OAI21X1_584 (.gnd(gnd), .A(_2131_), .Y(_902_), .vdd(vdd), .B(_2101__bF_buf0), .C(_2132_), );
  INVX2 INVX2_273 (.gnd(gnd), .A(regs_7__16_), .Y(_2133_), .vdd(vdd), );
  NAND2X1 NAND2X1_276 (.gnd(gnd), .A(wdata[16]), .Y(_2134_), .vdd(vdd), .B(_2101__bF_buf7), );
  OAI21X1 OAI21X1_585 (.gnd(gnd), .A(_2133_), .Y(_903_), .vdd(vdd), .B(_2101__bF_buf6), .C(_2134_), );
  INVX2 INVX2_274 (.gnd(gnd), .A(regs_7__17_), .Y(_2135_), .vdd(vdd), );
  NAND2X1 NAND2X1_277 (.gnd(gnd), .A(wdata[17]), .Y(_2136_), .vdd(vdd), .B(_2101__bF_buf5), );
  OAI21X1 OAI21X1_586 (.gnd(gnd), .A(_2135_), .Y(_904_), .vdd(vdd), .B(_2101__bF_buf4), .C(_2136_), );
  INVX2 INVX2_275 (.gnd(gnd), .A(regs_7__18_), .Y(_2137_), .vdd(vdd), );
  NAND2X1 NAND2X1_278 (.gnd(gnd), .A(wdata[18]), .Y(_2138_), .vdd(vdd), .B(_2101__bF_buf3), );
  OAI21X1 OAI21X1_587 (.gnd(gnd), .A(_2137_), .Y(_905_), .vdd(vdd), .B(_2101__bF_buf2), .C(_2138_), );
  INVX2 INVX2_276 (.gnd(gnd), .A(regs_7__19_), .Y(_2139_), .vdd(vdd), );
  NAND2X1 NAND2X1_279 (.gnd(gnd), .A(wdata[19]), .Y(_2140_), .vdd(vdd), .B(_2101__bF_buf1), );
  OAI21X1 OAI21X1_588 (.gnd(gnd), .A(_2139_), .Y(_906_), .vdd(vdd), .B(_2101__bF_buf0), .C(_2140_), );
  INVX2 INVX2_277 (.gnd(gnd), .A(regs_7__20_), .Y(_2141_), .vdd(vdd), );
  NAND2X1 NAND2X1_280 (.gnd(gnd), .A(wdata[20]), .Y(_2142_), .vdd(vdd), .B(_2101__bF_buf7), );
  OAI21X1 OAI21X1_589 (.gnd(gnd), .A(_2141_), .Y(_908_), .vdd(vdd), .B(_2101__bF_buf6), .C(_2142_), );
  INVX2 INVX2_278 (.gnd(gnd), .A(regs_7__21_), .Y(_2143_), .vdd(vdd), );
  NAND2X1 NAND2X1_281 (.gnd(gnd), .A(wdata[21]), .Y(_2144_), .vdd(vdd), .B(_2101__bF_buf5), );
  OAI21X1 OAI21X1_590 (.gnd(gnd), .A(_2143_), .Y(_909_), .vdd(vdd), .B(_2101__bF_buf4), .C(_2144_), );
  INVX2 INVX2_279 (.gnd(gnd), .A(regs_7__22_), .Y(_2145_), .vdd(vdd), );
  NAND2X1 NAND2X1_282 (.gnd(gnd), .A(wdata[22]), .Y(_2146_), .vdd(vdd), .B(_2101__bF_buf3), );
  OAI21X1 OAI21X1_591 (.gnd(gnd), .A(_2145_), .Y(_910_), .vdd(vdd), .B(_2101__bF_buf2), .C(_2146_), );
  INVX2 INVX2_280 (.gnd(gnd), .A(regs_7__23_), .Y(_2147_), .vdd(vdd), );
  NAND2X1 NAND2X1_283 (.gnd(gnd), .A(wdata[23]), .Y(_2148_), .vdd(vdd), .B(_2101__bF_buf1), );
  OAI21X1 OAI21X1_592 (.gnd(gnd), .A(_2147_), .Y(_911_), .vdd(vdd), .B(_2101__bF_buf0), .C(_2148_), );
  INVX2 INVX2_281 (.gnd(gnd), .A(regs_7__24_), .Y(_2149_), .vdd(vdd), );
  NAND2X1 NAND2X1_284 (.gnd(gnd), .A(wdata[24]), .Y(_2150_), .vdd(vdd), .B(_2101__bF_buf7), );
  OAI21X1 OAI21X1_593 (.gnd(gnd), .A(_2149_), .Y(_912_), .vdd(vdd), .B(_2101__bF_buf6), .C(_2150_), );
  INVX2 INVX2_282 (.gnd(gnd), .A(regs_7__25_), .Y(_2151_), .vdd(vdd), );
  NAND2X1 NAND2X1_285 (.gnd(gnd), .A(wdata[25]), .Y(_2152_), .vdd(vdd), .B(_2101__bF_buf5), );
  OAI21X1 OAI21X1_594 (.gnd(gnd), .A(_2151_), .Y(_913_), .vdd(vdd), .B(_2101__bF_buf4), .C(_2152_), );
  INVX2 INVX2_283 (.gnd(gnd), .A(regs_7__26_), .Y(_2153_), .vdd(vdd), );
  NAND2X1 NAND2X1_286 (.gnd(gnd), .A(wdata[26]), .Y(_2154_), .vdd(vdd), .B(_2101__bF_buf3), );
  OAI21X1 OAI21X1_595 (.gnd(gnd), .A(_2153_), .Y(_914_), .vdd(vdd), .B(_2101__bF_buf2), .C(_2154_), );
  INVX2 INVX2_284 (.gnd(gnd), .A(regs_7__27_), .Y(_2155_), .vdd(vdd), );
  NAND2X1 NAND2X1_287 (.gnd(gnd), .A(wdata[27]), .Y(_2156_), .vdd(vdd), .B(_2101__bF_buf1), );
  OAI21X1 OAI21X1_596 (.gnd(gnd), .A(_2155_), .Y(_915_), .vdd(vdd), .B(_2101__bF_buf0), .C(_2156_), );
  INVX2 INVX2_285 (.gnd(gnd), .A(regs_7__28_), .Y(_2157_), .vdd(vdd), );
  NAND2X1 NAND2X1_288 (.gnd(gnd), .A(wdata[28]), .Y(_2158_), .vdd(vdd), .B(_2101__bF_buf7), );
  OAI21X1 OAI21X1_597 (.gnd(gnd), .A(_2157_), .Y(_916_), .vdd(vdd), .B(_2101__bF_buf6), .C(_2158_), );
  INVX2 INVX2_286 (.gnd(gnd), .A(regs_7__29_), .Y(_2159_), .vdd(vdd), );
  NAND2X1 NAND2X1_289 (.gnd(gnd), .A(wdata[29]), .Y(_2160_), .vdd(vdd), .B(_2101__bF_buf5), );
  OAI21X1 OAI21X1_598 (.gnd(gnd), .A(_2159_), .Y(_917_), .vdd(vdd), .B(_2101__bF_buf4), .C(_2160_), );
  INVX2 INVX2_287 (.gnd(gnd), .A(regs_7__30_), .Y(_2161_), .vdd(vdd), );
  NAND2X1 NAND2X1_290 (.gnd(gnd), .A(wdata[30]), .Y(_2162_), .vdd(vdd), .B(_2101__bF_buf3), );
  OAI21X1 OAI21X1_599 (.gnd(gnd), .A(_2161_), .Y(_919_), .vdd(vdd), .B(_2101__bF_buf2), .C(_2162_), );
  INVX2 INVX2_288 (.gnd(gnd), .A(regs_7__31_), .Y(_2163_), .vdd(vdd), );
  NAND2X1 NAND2X1_291 (.gnd(gnd), .A(wdata[31]), .Y(_2164_), .vdd(vdd), .B(_2101__bF_buf1), );
  OAI21X1 OAI21X1_600 (.gnd(gnd), .A(_2163_), .Y(_920_), .vdd(vdd), .B(_2101__bF_buf0), .C(_2164_), );
  NAND2X1 NAND2X1_292 (.gnd(gnd), .A(_998_), .Y(_2165_), .vdd(vdd), .B(_2099_), );
  OAI21X1 OAI21X1_601 (.gnd(gnd), .A(_1001__bF_buf5), .Y(_2166_), .vdd(vdd), .B(_2100__bF_buf7), .C(regs_6__0_), );
  OAI21X1 OAI21X1_602 (.gnd(gnd), .A(_992__bF_buf3), .Y(_864_), .vdd(vdd), .B(_2165__bF_buf4), .C(_2166_), );
  OAI21X1 OAI21X1_603 (.gnd(gnd), .A(_1001__bF_buf4), .Y(_2167_), .vdd(vdd), .B(_2100__bF_buf6), .C(regs_6__1_), );
  OAI21X1 OAI21X1_604 (.gnd(gnd), .A(_1003__bF_buf3), .Y(_875_), .vdd(vdd), .B(_2165__bF_buf3), .C(_2167_), );
  OAI21X1 OAI21X1_605 (.gnd(gnd), .A(_1001__bF_buf3), .Y(_2168_), .vdd(vdd), .B(_2100__bF_buf5), .C(regs_6__2_), );
  OAI21X1 OAI21X1_606 (.gnd(gnd), .A(_1005__bF_buf3), .Y(_886_), .vdd(vdd), .B(_2165__bF_buf2), .C(_2168_), );
  OAI21X1 OAI21X1_607 (.gnd(gnd), .A(_1001__bF_buf2), .Y(_2169_), .vdd(vdd), .B(_2100__bF_buf4), .C(regs_6__3_), );
  OAI21X1 OAI21X1_608 (.gnd(gnd), .A(_1007__bF_buf3), .Y(_889_), .vdd(vdd), .B(_2165__bF_buf1), .C(_2169_), );
  OAI21X1 OAI21X1_609 (.gnd(gnd), .A(_1001__bF_buf1), .Y(_2170_), .vdd(vdd), .B(_2100__bF_buf3), .C(regs_6__4_), );
  OAI21X1 OAI21X1_610 (.gnd(gnd), .A(_1009__bF_buf2), .Y(_890_), .vdd(vdd), .B(_2165__bF_buf0), .C(_2170_), );
  OAI21X1 OAI21X1_611 (.gnd(gnd), .A(_1001__bF_buf0), .Y(_2171_), .vdd(vdd), .B(_2100__bF_buf2), .C(regs_6__5_), );
  OAI21X1 OAI21X1_612 (.gnd(gnd), .A(_1011__bF_buf2), .Y(_891_), .vdd(vdd), .B(_2165__bF_buf4), .C(_2171_), );
  OAI21X1 OAI21X1_613 (.gnd(gnd), .A(_1001__bF_buf9), .Y(_2172_), .vdd(vdd), .B(_2100__bF_buf1), .C(regs_6__6_), );
  OAI21X1 OAI21X1_614 (.gnd(gnd), .A(_1013__bF_buf2), .Y(_892_), .vdd(vdd), .B(_2165__bF_buf3), .C(_2172_), );
  OAI21X1 OAI21X1_615 (.gnd(gnd), .A(_1001__bF_buf8), .Y(_2173_), .vdd(vdd), .B(_2100__bF_buf0), .C(regs_6__7_), );
  OAI21X1 OAI21X1_616 (.gnd(gnd), .A(_1015__bF_buf2), .Y(_893_), .vdd(vdd), .B(_2165__bF_buf2), .C(_2173_), );
  OAI21X1 OAI21X1_617 (.gnd(gnd), .A(_1001__bF_buf7), .Y(_2174_), .vdd(vdd), .B(_2100__bF_buf8), .C(regs_6__8_), );
  OAI21X1 OAI21X1_618 (.gnd(gnd), .A(_1017__bF_buf2), .Y(_894_), .vdd(vdd), .B(_2165__bF_buf1), .C(_2174_), );
  OAI21X1 OAI21X1_619 (.gnd(gnd), .A(_1001__bF_buf6), .Y(_2175_), .vdd(vdd), .B(_2100__bF_buf7), .C(regs_6__9_), );
  OAI21X1 OAI21X1_620 (.gnd(gnd), .A(_1019__bF_buf2), .Y(_895_), .vdd(vdd), .B(_2165__bF_buf0), .C(_2175_), );
  OAI21X1 OAI21X1_621 (.gnd(gnd), .A(_1001__bF_buf5), .Y(_2176_), .vdd(vdd), .B(_2100__bF_buf6), .C(regs_6__10_), );
  OAI21X1 OAI21X1_622 (.gnd(gnd), .A(_1021__bF_buf2), .Y(_865_), .vdd(vdd), .B(_2165__bF_buf4), .C(_2176_), );
  OAI21X1 OAI21X1_623 (.gnd(gnd), .A(_1001__bF_buf4), .Y(_2177_), .vdd(vdd), .B(_2100__bF_buf5), .C(regs_6__11_), );
  OAI21X1 OAI21X1_624 (.gnd(gnd), .A(_1023__bF_buf2), .Y(_866_), .vdd(vdd), .B(_2165__bF_buf3), .C(_2177_), );
  OAI21X1 OAI21X1_625 (.gnd(gnd), .A(_1001__bF_buf3), .Y(_2178_), .vdd(vdd), .B(_2100__bF_buf4), .C(regs_6__12_), );
  OAI21X1 OAI21X1_626 (.gnd(gnd), .A(_1025__bF_buf2), .Y(_867_), .vdd(vdd), .B(_2165__bF_buf2), .C(_2178_), );
  OAI21X1 OAI21X1_627 (.gnd(gnd), .A(_1001__bF_buf2), .Y(_2179_), .vdd(vdd), .B(_2100__bF_buf3), .C(regs_6__13_), );
  OAI21X1 OAI21X1_628 (.gnd(gnd), .A(_1027__bF_buf2), .Y(_868_), .vdd(vdd), .B(_2165__bF_buf1), .C(_2179_), );
  OAI21X1 OAI21X1_629 (.gnd(gnd), .A(_1001__bF_buf1), .Y(_2180_), .vdd(vdd), .B(_2100__bF_buf2), .C(regs_6__14_), );
  OAI21X1 OAI21X1_630 (.gnd(gnd), .A(_1029__bF_buf2), .Y(_869_), .vdd(vdd), .B(_2165__bF_buf0), .C(_2180_), );
  OAI21X1 OAI21X1_631 (.gnd(gnd), .A(_1001__bF_buf0), .Y(_2181_), .vdd(vdd), .B(_2100__bF_buf1), .C(regs_6__15_), );
  OAI21X1 OAI21X1_632 (.gnd(gnd), .A(_1031__bF_buf2), .Y(_870_), .vdd(vdd), .B(_2165__bF_buf4), .C(_2181_), );
  OAI21X1 OAI21X1_633 (.gnd(gnd), .A(_1001__bF_buf9), .Y(_2182_), .vdd(vdd), .B(_2100__bF_buf0), .C(regs_6__16_), );
  OAI21X1 OAI21X1_634 (.gnd(gnd), .A(_1033__bF_buf2), .Y(_871_), .vdd(vdd), .B(_2165__bF_buf3), .C(_2182_), );
  OAI21X1 OAI21X1_635 (.gnd(gnd), .A(_1001__bF_buf8), .Y(_2183_), .vdd(vdd), .B(_2100__bF_buf8), .C(regs_6__17_), );
  OAI21X1 OAI21X1_636 (.gnd(gnd), .A(_1035__bF_buf2), .Y(_872_), .vdd(vdd), .B(_2165__bF_buf2), .C(_2183_), );
  OAI21X1 OAI21X1_637 (.gnd(gnd), .A(_1001__bF_buf7), .Y(_2184_), .vdd(vdd), .B(_2100__bF_buf7), .C(regs_6__18_), );
  OAI21X1 OAI21X1_638 (.gnd(gnd), .A(_1037__bF_buf2), .Y(_873_), .vdd(vdd), .B(_2165__bF_buf1), .C(_2184_), );
  OAI21X1 OAI21X1_639 (.gnd(gnd), .A(_1001__bF_buf6), .Y(_2185_), .vdd(vdd), .B(_2100__bF_buf6), .C(regs_6__19_), );
  OAI21X1 OAI21X1_640 (.gnd(gnd), .A(_1039__bF_buf2), .Y(_874_), .vdd(vdd), .B(_2165__bF_buf0), .C(_2185_), );
  OAI21X1 OAI21X1_641 (.gnd(gnd), .A(_1001__bF_buf5), .Y(_2186_), .vdd(vdd), .B(_2100__bF_buf5), .C(regs_6__20_), );
  OAI21X1 OAI21X1_642 (.gnd(gnd), .A(_1041__bF_buf2), .Y(_876_), .vdd(vdd), .B(_2165__bF_buf4), .C(_2186_), );
  OAI21X1 OAI21X1_643 (.gnd(gnd), .A(_1001__bF_buf4), .Y(_2187_), .vdd(vdd), .B(_2100__bF_buf4), .C(regs_6__21_), );
  OAI21X1 OAI21X1_644 (.gnd(gnd), .A(_1043__bF_buf2), .Y(_877_), .vdd(vdd), .B(_2165__bF_buf3), .C(_2187_), );
  OAI21X1 OAI21X1_645 (.gnd(gnd), .A(_1001__bF_buf3), .Y(_2188_), .vdd(vdd), .B(_2100__bF_buf3), .C(regs_6__22_), );
  OAI21X1 OAI21X1_646 (.gnd(gnd), .A(_1045__bF_buf2), .Y(_878_), .vdd(vdd), .B(_2165__bF_buf2), .C(_2188_), );
  OAI21X1 OAI21X1_647 (.gnd(gnd), .A(_1001__bF_buf2), .Y(_2189_), .vdd(vdd), .B(_2100__bF_buf2), .C(regs_6__23_), );
  OAI21X1 OAI21X1_648 (.gnd(gnd), .A(_1047__bF_buf2), .Y(_879_), .vdd(vdd), .B(_2165__bF_buf1), .C(_2189_), );
  OAI21X1 OAI21X1_649 (.gnd(gnd), .A(_1001__bF_buf1), .Y(_2190_), .vdd(vdd), .B(_2100__bF_buf1), .C(regs_6__24_), );
  OAI21X1 OAI21X1_650 (.gnd(gnd), .A(_1049__bF_buf2), .Y(_880_), .vdd(vdd), .B(_2165__bF_buf0), .C(_2190_), );
  OAI21X1 OAI21X1_651 (.gnd(gnd), .A(_1001__bF_buf0), .Y(_2191_), .vdd(vdd), .B(_2100__bF_buf0), .C(regs_6__25_), );
  OAI21X1 OAI21X1_652 (.gnd(gnd), .A(_1051__bF_buf2), .Y(_881_), .vdd(vdd), .B(_2165__bF_buf4), .C(_2191_), );
  OAI21X1 OAI21X1_653 (.gnd(gnd), .A(_1001__bF_buf9), .Y(_2192_), .vdd(vdd), .B(_2100__bF_buf8), .C(regs_6__26_), );
  OAI21X1 OAI21X1_654 (.gnd(gnd), .A(_1053__bF_buf2), .Y(_882_), .vdd(vdd), .B(_2165__bF_buf3), .C(_2192_), );
  OAI21X1 OAI21X1_655 (.gnd(gnd), .A(_1001__bF_buf8), .Y(_2193_), .vdd(vdd), .B(_2100__bF_buf7), .C(regs_6__27_), );
  OAI21X1 OAI21X1_656 (.gnd(gnd), .A(_1055__bF_buf2), .Y(_883_), .vdd(vdd), .B(_2165__bF_buf2), .C(_2193_), );
  OAI21X1 OAI21X1_657 (.gnd(gnd), .A(_1001__bF_buf7), .Y(_2194_), .vdd(vdd), .B(_2100__bF_buf6), .C(regs_6__28_), );
  OAI21X1 OAI21X1_658 (.gnd(gnd), .A(_1057__bF_buf2), .Y(_884_), .vdd(vdd), .B(_2165__bF_buf1), .C(_2194_), );
  OAI21X1 OAI21X1_659 (.gnd(gnd), .A(_1001__bF_buf6), .Y(_2195_), .vdd(vdd), .B(_2100__bF_buf5), .C(regs_6__29_), );
  OAI21X1 OAI21X1_660 (.gnd(gnd), .A(_1059__bF_buf2), .Y(_885_), .vdd(vdd), .B(_2165__bF_buf0), .C(_2195_), );
  OAI21X1 OAI21X1_661 (.gnd(gnd), .A(_1001__bF_buf5), .Y(_2196_), .vdd(vdd), .B(_2100__bF_buf4), .C(regs_6__30_), );
  OAI21X1 OAI21X1_662 (.gnd(gnd), .A(_1061__bF_buf2), .Y(_887_), .vdd(vdd), .B(_2165__bF_buf4), .C(_2196_), );
  OAI21X1 OAI21X1_663 (.gnd(gnd), .A(_1001__bF_buf4), .Y(_2197_), .vdd(vdd), .B(_2100__bF_buf3), .C(regs_6__31_), );
  OAI21X1 OAI21X1_664 (.gnd(gnd), .A(_1063__bF_buf2), .Y(_888_), .vdd(vdd), .B(_2165__bF_buf3), .C(_2197_), );
  NAND2X1 NAND2X1_293 (.gnd(gnd), .A(_2099_), .Y(_2198_), .vdd(vdd), .B(_1068_), );
  OAI21X1 OAI21X1_665 (.gnd(gnd), .A(_1070__bF_buf6), .Y(_2199_), .vdd(vdd), .B(_2100__bF_buf2), .C(regs_5__0_), );
  OAI21X1 OAI21X1_666 (.gnd(gnd), .A(_992__bF_buf2), .Y(_832_), .vdd(vdd), .B(_2198__bF_buf4), .C(_2199_), );
  OAI21X1 OAI21X1_667 (.gnd(gnd), .A(_1070__bF_buf5), .Y(_2200_), .vdd(vdd), .B(_2100__bF_buf1), .C(regs_5__1_), );
  OAI21X1 OAI21X1_668 (.gnd(gnd), .A(_1003__bF_buf2), .Y(_843_), .vdd(vdd), .B(_2198__bF_buf3), .C(_2200_), );
  OAI21X1 OAI21X1_669 (.gnd(gnd), .A(_1070__bF_buf4), .Y(_2201_), .vdd(vdd), .B(_2100__bF_buf0), .C(regs_5__2_), );
  OAI21X1 OAI21X1_670 (.gnd(gnd), .A(_1005__bF_buf2), .Y(_854_), .vdd(vdd), .B(_2198__bF_buf2), .C(_2201_), );
  OAI21X1 OAI21X1_671 (.gnd(gnd), .A(_1070__bF_buf3), .Y(_2202_), .vdd(vdd), .B(_2100__bF_buf8), .C(regs_5__3_), );
  OAI21X1 OAI21X1_672 (.gnd(gnd), .A(_1007__bF_buf2), .Y(_857_), .vdd(vdd), .B(_2198__bF_buf1), .C(_2202_), );
  OAI21X1 OAI21X1_673 (.gnd(gnd), .A(_1070__bF_buf2), .Y(_2203_), .vdd(vdd), .B(_2100__bF_buf7), .C(regs_5__4_), );
  OAI21X1 OAI21X1_674 (.gnd(gnd), .A(_1009__bF_buf1), .Y(_858_), .vdd(vdd), .B(_2198__bF_buf0), .C(_2203_), );
  OAI21X1 OAI21X1_675 (.gnd(gnd), .A(_1070__bF_buf1), .Y(_2204_), .vdd(vdd), .B(_2100__bF_buf6), .C(regs_5__5_), );
  OAI21X1 OAI21X1_676 (.gnd(gnd), .A(_1011__bF_buf1), .Y(_859_), .vdd(vdd), .B(_2198__bF_buf4), .C(_2204_), );
  OAI21X1 OAI21X1_677 (.gnd(gnd), .A(_1070__bF_buf0), .Y(_2205_), .vdd(vdd), .B(_2100__bF_buf5), .C(regs_5__6_), );
  OAI21X1 OAI21X1_678 (.gnd(gnd), .A(_1013__bF_buf1), .Y(_860_), .vdd(vdd), .B(_2198__bF_buf3), .C(_2205_), );
  OAI21X1 OAI21X1_679 (.gnd(gnd), .A(_1070__bF_buf10), .Y(_2206_), .vdd(vdd), .B(_2100__bF_buf4), .C(regs_5__7_), );
  OAI21X1 OAI21X1_680 (.gnd(gnd), .A(_1015__bF_buf1), .Y(_861_), .vdd(vdd), .B(_2198__bF_buf2), .C(_2206_), );
  OAI21X1 OAI21X1_681 (.gnd(gnd), .A(_1070__bF_buf9), .Y(_2207_), .vdd(vdd), .B(_2100__bF_buf3), .C(regs_5__8_), );
  OAI21X1 OAI21X1_682 (.gnd(gnd), .A(_1017__bF_buf1), .Y(_862_), .vdd(vdd), .B(_2198__bF_buf1), .C(_2207_), );
  OAI21X1 OAI21X1_683 (.gnd(gnd), .A(_1070__bF_buf8), .Y(_2208_), .vdd(vdd), .B(_2100__bF_buf2), .C(regs_5__9_), );
  OAI21X1 OAI21X1_684 (.gnd(gnd), .A(_1019__bF_buf1), .Y(_863_), .vdd(vdd), .B(_2198__bF_buf0), .C(_2208_), );
  OAI21X1 OAI21X1_685 (.gnd(gnd), .A(_1070__bF_buf7), .Y(_2209_), .vdd(vdd), .B(_2100__bF_buf1), .C(regs_5__10_), );
  OAI21X1 OAI21X1_686 (.gnd(gnd), .A(_1021__bF_buf1), .Y(_833_), .vdd(vdd), .B(_2198__bF_buf4), .C(_2209_), );
  OAI21X1 OAI21X1_687 (.gnd(gnd), .A(_1070__bF_buf6), .Y(_2210_), .vdd(vdd), .B(_2100__bF_buf0), .C(regs_5__11_), );
  OAI21X1 OAI21X1_688 (.gnd(gnd), .A(_1023__bF_buf1), .Y(_834_), .vdd(vdd), .B(_2198__bF_buf3), .C(_2210_), );
  OAI21X1 OAI21X1_689 (.gnd(gnd), .A(_1070__bF_buf5), .Y(_2211_), .vdd(vdd), .B(_2100__bF_buf8), .C(regs_5__12_), );
  OAI21X1 OAI21X1_690 (.gnd(gnd), .A(_1025__bF_buf1), .Y(_835_), .vdd(vdd), .B(_2198__bF_buf2), .C(_2211_), );
  OAI21X1 OAI21X1_691 (.gnd(gnd), .A(_1070__bF_buf4), .Y(_2212_), .vdd(vdd), .B(_2100__bF_buf7), .C(regs_5__13_), );
  OAI21X1 OAI21X1_692 (.gnd(gnd), .A(_1027__bF_buf1), .Y(_836_), .vdd(vdd), .B(_2198__bF_buf1), .C(_2212_), );
  OAI21X1 OAI21X1_693 (.gnd(gnd), .A(_1070__bF_buf3), .Y(_2213_), .vdd(vdd), .B(_2100__bF_buf6), .C(regs_5__14_), );
  OAI21X1 OAI21X1_694 (.gnd(gnd), .A(_1029__bF_buf1), .Y(_837_), .vdd(vdd), .B(_2198__bF_buf0), .C(_2213_), );
  OAI21X1 OAI21X1_695 (.gnd(gnd), .A(_1070__bF_buf2), .Y(_2214_), .vdd(vdd), .B(_2100__bF_buf5), .C(regs_5__15_), );
  OAI21X1 OAI21X1_696 (.gnd(gnd), .A(_1031__bF_buf1), .Y(_838_), .vdd(vdd), .B(_2198__bF_buf4), .C(_2214_), );
  OAI21X1 OAI21X1_697 (.gnd(gnd), .A(_1070__bF_buf1), .Y(_2215_), .vdd(vdd), .B(_2100__bF_buf4), .C(regs_5__16_), );
  OAI21X1 OAI21X1_698 (.gnd(gnd), .A(_1033__bF_buf1), .Y(_839_), .vdd(vdd), .B(_2198__bF_buf3), .C(_2215_), );
  OAI21X1 OAI21X1_699 (.gnd(gnd), .A(_1070__bF_buf0), .Y(_2216_), .vdd(vdd), .B(_2100__bF_buf3), .C(regs_5__17_), );
  OAI21X1 OAI21X1_700 (.gnd(gnd), .A(_1035__bF_buf1), .Y(_840_), .vdd(vdd), .B(_2198__bF_buf2), .C(_2216_), );
  OAI21X1 OAI21X1_701 (.gnd(gnd), .A(_1070__bF_buf10), .Y(_2217_), .vdd(vdd), .B(_2100__bF_buf2), .C(regs_5__18_), );
  OAI21X1 OAI21X1_702 (.gnd(gnd), .A(_1037__bF_buf1), .Y(_841_), .vdd(vdd), .B(_2198__bF_buf1), .C(_2217_), );
  OAI21X1 OAI21X1_703 (.gnd(gnd), .A(_1070__bF_buf9), .Y(_2218_), .vdd(vdd), .B(_2100__bF_buf1), .C(regs_5__19_), );
  OAI21X1 OAI21X1_704 (.gnd(gnd), .A(_1039__bF_buf1), .Y(_842_), .vdd(vdd), .B(_2198__bF_buf0), .C(_2218_), );
  OAI21X1 OAI21X1_705 (.gnd(gnd), .A(_1070__bF_buf8), .Y(_2219_), .vdd(vdd), .B(_2100__bF_buf0), .C(regs_5__20_), );
  OAI21X1 OAI21X1_706 (.gnd(gnd), .A(_1041__bF_buf1), .Y(_844_), .vdd(vdd), .B(_2198__bF_buf4), .C(_2219_), );
  OAI21X1 OAI21X1_707 (.gnd(gnd), .A(_1070__bF_buf7), .Y(_2220_), .vdd(vdd), .B(_2100__bF_buf8), .C(regs_5__21_), );
  OAI21X1 OAI21X1_708 (.gnd(gnd), .A(_1043__bF_buf1), .Y(_845_), .vdd(vdd), .B(_2198__bF_buf3), .C(_2220_), );
  OAI21X1 OAI21X1_709 (.gnd(gnd), .A(_1070__bF_buf6), .Y(_2221_), .vdd(vdd), .B(_2100__bF_buf7), .C(regs_5__22_), );
  OAI21X1 OAI21X1_710 (.gnd(gnd), .A(_1045__bF_buf1), .Y(_846_), .vdd(vdd), .B(_2198__bF_buf2), .C(_2221_), );
  OAI21X1 OAI21X1_711 (.gnd(gnd), .A(_1070__bF_buf5), .Y(_2222_), .vdd(vdd), .B(_2100__bF_buf6), .C(regs_5__23_), );
  OAI21X1 OAI21X1_712 (.gnd(gnd), .A(_1047__bF_buf1), .Y(_847_), .vdd(vdd), .B(_2198__bF_buf1), .C(_2222_), );
  OAI21X1 OAI21X1_713 (.gnd(gnd), .A(_1070__bF_buf4), .Y(_2223_), .vdd(vdd), .B(_2100__bF_buf5), .C(regs_5__24_), );
  OAI21X1 OAI21X1_714 (.gnd(gnd), .A(_1049__bF_buf1), .Y(_848_), .vdd(vdd), .B(_2198__bF_buf0), .C(_2223_), );
  OAI21X1 OAI21X1_715 (.gnd(gnd), .A(_1070__bF_buf3), .Y(_2224_), .vdd(vdd), .B(_2100__bF_buf4), .C(regs_5__25_), );
  OAI21X1 OAI21X1_716 (.gnd(gnd), .A(_1051__bF_buf1), .Y(_849_), .vdd(vdd), .B(_2198__bF_buf4), .C(_2224_), );
  OAI21X1 OAI21X1_717 (.gnd(gnd), .A(_1070__bF_buf2), .Y(_2225_), .vdd(vdd), .B(_2100__bF_buf3), .C(regs_5__26_), );
  OAI21X1 OAI21X1_718 (.gnd(gnd), .A(_1053__bF_buf1), .Y(_850_), .vdd(vdd), .B(_2198__bF_buf3), .C(_2225_), );
  OAI21X1 OAI21X1_719 (.gnd(gnd), .A(_1070__bF_buf1), .Y(_2226_), .vdd(vdd), .B(_2100__bF_buf2), .C(regs_5__27_), );
  OAI21X1 OAI21X1_720 (.gnd(gnd), .A(_1055__bF_buf1), .Y(_851_), .vdd(vdd), .B(_2198__bF_buf2), .C(_2226_), );
  OAI21X1 OAI21X1_721 (.gnd(gnd), .A(_1070__bF_buf0), .Y(_2227_), .vdd(vdd), .B(_2100__bF_buf1), .C(regs_5__28_), );
  OAI21X1 OAI21X1_722 (.gnd(gnd), .A(_1057__bF_buf1), .Y(_852_), .vdd(vdd), .B(_2198__bF_buf1), .C(_2227_), );
  OAI21X1 OAI21X1_723 (.gnd(gnd), .A(_1070__bF_buf10), .Y(_2228_), .vdd(vdd), .B(_2100__bF_buf0), .C(regs_5__29_), );
  OAI21X1 OAI21X1_724 (.gnd(gnd), .A(_1059__bF_buf1), .Y(_853_), .vdd(vdd), .B(_2198__bF_buf0), .C(_2228_), );
  OAI21X1 OAI21X1_725 (.gnd(gnd), .A(_1070__bF_buf9), .Y(_2229_), .vdd(vdd), .B(_2100__bF_buf8), .C(regs_5__30_), );
  OAI21X1 OAI21X1_726 (.gnd(gnd), .A(_1061__bF_buf1), .Y(_855_), .vdd(vdd), .B(_2198__bF_buf4), .C(_2229_), );
  OAI21X1 OAI21X1_727 (.gnd(gnd), .A(_1070__bF_buf8), .Y(_2230_), .vdd(vdd), .B(_2100__bF_buf7), .C(regs_5__31_), );
  OAI21X1 OAI21X1_728 (.gnd(gnd), .A(_1063__bF_buf1), .Y(_856_), .vdd(vdd), .B(_2198__bF_buf3), .C(_2230_), );
  NAND2X1 NAND2X1_294 (.gnd(gnd), .A(_2099_), .Y(_2231_), .vdd(vdd), .B(_1273_), );
  OAI21X1 OAI21X1_729 (.gnd(gnd), .A(_2100__bF_buf6), .Y(_2232_), .vdd(vdd), .B(_1104__bF_buf4), .C(regs_4__0_), );
  OAI21X1 OAI21X1_730 (.gnd(gnd), .A(_2231__bF_buf4), .Y(_800_), .vdd(vdd), .B(_992__bF_buf1), .C(_2232_), );
  OAI21X1 OAI21X1_731 (.gnd(gnd), .A(_2100__bF_buf5), .Y(_2233_), .vdd(vdd), .B(_1104__bF_buf3), .C(regs_4__1_), );
  OAI21X1 OAI21X1_732 (.gnd(gnd), .A(_2231__bF_buf3), .Y(_811_), .vdd(vdd), .B(_1003__bF_buf1), .C(_2233_), );
  OAI21X1 OAI21X1_733 (.gnd(gnd), .A(_2100__bF_buf4), .Y(_2234_), .vdd(vdd), .B(_1104__bF_buf2), .C(regs_4__2_), );
  OAI21X1 OAI21X1_734 (.gnd(gnd), .A(_2231__bF_buf2), .Y(_822_), .vdd(vdd), .B(_1005__bF_buf1), .C(_2234_), );
  OAI21X1 OAI21X1_735 (.gnd(gnd), .A(_2100__bF_buf3), .Y(_2235_), .vdd(vdd), .B(_1104__bF_buf1), .C(regs_4__3_), );
  OAI21X1 OAI21X1_736 (.gnd(gnd), .A(_2231__bF_buf1), .Y(_825_), .vdd(vdd), .B(_1007__bF_buf1), .C(_2235_), );
  OAI21X1 OAI21X1_737 (.gnd(gnd), .A(_2100__bF_buf2), .Y(_2236_), .vdd(vdd), .B(_1104__bF_buf0), .C(regs_4__4_), );
  OAI21X1 OAI21X1_738 (.gnd(gnd), .A(_2231__bF_buf0), .Y(_826_), .vdd(vdd), .B(_1009__bF_buf0), .C(_2236_), );
  OAI21X1 OAI21X1_739 (.gnd(gnd), .A(_2100__bF_buf1), .Y(_2237_), .vdd(vdd), .B(_1104__bF_buf14), .C(regs_4__5_), );
  OAI21X1 OAI21X1_740 (.gnd(gnd), .A(_2231__bF_buf4), .Y(_827_), .vdd(vdd), .B(_1011__bF_buf0), .C(_2237_), );
  OAI21X1 OAI21X1_741 (.gnd(gnd), .A(_2100__bF_buf0), .Y(_2238_), .vdd(vdd), .B(_1104__bF_buf13), .C(regs_4__6_), );
  OAI21X1 OAI21X1_742 (.gnd(gnd), .A(_2231__bF_buf3), .Y(_828_), .vdd(vdd), .B(_1013__bF_buf0), .C(_2238_), );
  OAI21X1 OAI21X1_743 (.gnd(gnd), .A(_2100__bF_buf8), .Y(_2239_), .vdd(vdd), .B(_1104__bF_buf12), .C(regs_4__7_), );
  OAI21X1 OAI21X1_744 (.gnd(gnd), .A(_2231__bF_buf2), .Y(_829_), .vdd(vdd), .B(_1015__bF_buf0), .C(_2239_), );
  OAI21X1 OAI21X1_745 (.gnd(gnd), .A(_2100__bF_buf7), .Y(_2240_), .vdd(vdd), .B(_1104__bF_buf11), .C(regs_4__8_), );
  OAI21X1 OAI21X1_746 (.gnd(gnd), .A(_2231__bF_buf1), .Y(_830_), .vdd(vdd), .B(_1017__bF_buf0), .C(_2240_), );
  OAI21X1 OAI21X1_747 (.gnd(gnd), .A(_2100__bF_buf6), .Y(_2241_), .vdd(vdd), .B(_1104__bF_buf10), .C(regs_4__9_), );
  OAI21X1 OAI21X1_748 (.gnd(gnd), .A(_2231__bF_buf0), .Y(_831_), .vdd(vdd), .B(_1019__bF_buf0), .C(_2241_), );
  OAI21X1 OAI21X1_749 (.gnd(gnd), .A(_2100__bF_buf5), .Y(_2242_), .vdd(vdd), .B(_1104__bF_buf9), .C(regs_4__10_), );
  OAI21X1 OAI21X1_750 (.gnd(gnd), .A(_2231__bF_buf4), .Y(_801_), .vdd(vdd), .B(_1021__bF_buf0), .C(_2242_), );
  OAI21X1 OAI21X1_751 (.gnd(gnd), .A(_2100__bF_buf4), .Y(_2243_), .vdd(vdd), .B(_1104__bF_buf8), .C(regs_4__11_), );
  OAI21X1 OAI21X1_752 (.gnd(gnd), .A(_2231__bF_buf3), .Y(_802_), .vdd(vdd), .B(_1023__bF_buf0), .C(_2243_), );
  OAI21X1 OAI21X1_753 (.gnd(gnd), .A(_2100__bF_buf3), .Y(_2244_), .vdd(vdd), .B(_1104__bF_buf7), .C(regs_4__12_), );
  OAI21X1 OAI21X1_754 (.gnd(gnd), .A(_2231__bF_buf2), .Y(_803_), .vdd(vdd), .B(_1025__bF_buf0), .C(_2244_), );
  OAI21X1 OAI21X1_755 (.gnd(gnd), .A(_2100__bF_buf2), .Y(_2245_), .vdd(vdd), .B(_1104__bF_buf6), .C(regs_4__13_), );
  OAI21X1 OAI21X1_756 (.gnd(gnd), .A(_2231__bF_buf1), .Y(_804_), .vdd(vdd), .B(_1027__bF_buf0), .C(_2245_), );
  OAI21X1 OAI21X1_757 (.gnd(gnd), .A(_2100__bF_buf1), .Y(_2246_), .vdd(vdd), .B(_1104__bF_buf5), .C(regs_4__14_), );
  OAI21X1 OAI21X1_758 (.gnd(gnd), .A(_2231__bF_buf0), .Y(_805_), .vdd(vdd), .B(_1029__bF_buf0), .C(_2246_), );
  OAI21X1 OAI21X1_759 (.gnd(gnd), .A(_2100__bF_buf0), .Y(_2247_), .vdd(vdd), .B(_1104__bF_buf4), .C(regs_4__15_), );
  OAI21X1 OAI21X1_760 (.gnd(gnd), .A(_2231__bF_buf4), .Y(_806_), .vdd(vdd), .B(_1031__bF_buf0), .C(_2247_), );
  OAI21X1 OAI21X1_761 (.gnd(gnd), .A(_2100__bF_buf8), .Y(_2248_), .vdd(vdd), .B(_1104__bF_buf3), .C(regs_4__16_), );
  OAI21X1 OAI21X1_762 (.gnd(gnd), .A(_2231__bF_buf3), .Y(_807_), .vdd(vdd), .B(_1033__bF_buf0), .C(_2248_), );
  OAI21X1 OAI21X1_763 (.gnd(gnd), .A(_2100__bF_buf7), .Y(_2249_), .vdd(vdd), .B(_1104__bF_buf2), .C(regs_4__17_), );
  OAI21X1 OAI21X1_764 (.gnd(gnd), .A(_2231__bF_buf2), .Y(_808_), .vdd(vdd), .B(_1035__bF_buf0), .C(_2249_), );
  OAI21X1 OAI21X1_765 (.gnd(gnd), .A(_2100__bF_buf6), .Y(_2250_), .vdd(vdd), .B(_1104__bF_buf1), .C(regs_4__18_), );
  OAI21X1 OAI21X1_766 (.gnd(gnd), .A(_2231__bF_buf1), .Y(_809_), .vdd(vdd), .B(_1037__bF_buf0), .C(_2250_), );
  OAI21X1 OAI21X1_767 (.gnd(gnd), .A(_2100__bF_buf5), .Y(_2251_), .vdd(vdd), .B(_1104__bF_buf0), .C(regs_4__19_), );
  OAI21X1 OAI21X1_768 (.gnd(gnd), .A(_2231__bF_buf0), .Y(_810_), .vdd(vdd), .B(_1039__bF_buf0), .C(_2251_), );
  OAI21X1 OAI21X1_769 (.gnd(gnd), .A(_2100__bF_buf4), .Y(_2252_), .vdd(vdd), .B(_1104__bF_buf14), .C(regs_4__20_), );
  OAI21X1 OAI21X1_770 (.gnd(gnd), .A(_2231__bF_buf4), .Y(_812_), .vdd(vdd), .B(_1041__bF_buf0), .C(_2252_), );
  OAI21X1 OAI21X1_771 (.gnd(gnd), .A(_2100__bF_buf3), .Y(_2253_), .vdd(vdd), .B(_1104__bF_buf13), .C(regs_4__21_), );
  OAI21X1 OAI21X1_772 (.gnd(gnd), .A(_2231__bF_buf3), .Y(_813_), .vdd(vdd), .B(_1043__bF_buf0), .C(_2253_), );
  OAI21X1 OAI21X1_773 (.gnd(gnd), .A(_2100__bF_buf2), .Y(_2254_), .vdd(vdd), .B(_1104__bF_buf12), .C(regs_4__22_), );
  OAI21X1 OAI21X1_774 (.gnd(gnd), .A(_2231__bF_buf2), .Y(_814_), .vdd(vdd), .B(_1045__bF_buf0), .C(_2254_), );
  OAI21X1 OAI21X1_775 (.gnd(gnd), .A(_2100__bF_buf1), .Y(_2255_), .vdd(vdd), .B(_1104__bF_buf11), .C(regs_4__23_), );
  OAI21X1 OAI21X1_776 (.gnd(gnd), .A(_2231__bF_buf1), .Y(_815_), .vdd(vdd), .B(_1047__bF_buf0), .C(_2255_), );
  OAI21X1 OAI21X1_777 (.gnd(gnd), .A(_2100__bF_buf0), .Y(_2256_), .vdd(vdd), .B(_1104__bF_buf10), .C(regs_4__24_), );
  OAI21X1 OAI21X1_778 (.Y(_816_), .A(_2231__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1049__bF_buf0), .C(_2256_), );
  OAI21X1 OAI21X1_779 (.Y(_2257_), .A(_2100__bF_buf8), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf9), .C(regs_4__25_), );
  OAI21X1 OAI21X1_780 (.Y(_817_), .A(_2231__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1051__bF_buf0), .C(_2257_), );
  OAI21X1 OAI21X1_781 (.Y(_2258_), .A(_2100__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf8), .C(regs_4__26_), );
  OAI21X1 OAI21X1_782 (.Y(_818_), .A(_2231__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1053__bF_buf0), .C(_2258_), );
  OAI21X1 OAI21X1_783 (.Y(_2259_), .A(_2100__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf7), .C(regs_4__27_), );
  OAI21X1 OAI21X1_784 (.Y(_819_), .A(_2231__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1055__bF_buf0), .C(_2259_), );
  OAI21X1 OAI21X1_785 (.Y(_2260_), .A(_2100__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf6), .C(regs_4__28_), );
  OAI21X1 OAI21X1_786 (.Y(_820_), .A(_2231__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1057__bF_buf0), .C(_2260_), );
  OAI21X1 OAI21X1_787 (.Y(_2261_), .A(_2100__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf5), .C(regs_4__29_), );
  OAI21X1 OAI21X1_788 (.Y(_821_), .A(_2231__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1059__bF_buf0), .C(_2261_), );
  OAI21X1 OAI21X1_789 (.Y(_2262_), .A(_2100__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf4), .C(regs_4__30_), );
  OAI21X1 OAI21X1_790 (.Y(_823_), .A(_2231__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1061__bF_buf0), .C(_2262_), );
  OAI21X1 OAI21X1_791 (.Y(_2263_), .A(_2100__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1104__bF_buf3), .C(regs_4__31_), );
  OAI21X1 OAI21X1_792 (.Y(_824_), .A(_2231__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1063__bF_buf0), .C(_2263_), );
  OR2X2 OR2X2_9 (.Y(_2264_), .A(_2098_), .gnd(gnd), .vdd(vdd), .B(_1139_), );
  OR2X2 OR2X2_10 (.Y(_2265_), .A(_2264__bF_buf10), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf0), );
  OAI21X1 OAI21X1_793 (.Y(_2266_), .A(_2264__bF_buf9), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf5), .C(regs_3__0_), );
  OAI21X1 OAI21X1_794 (.Y(_768_), .A(_2265__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_992__bF_buf0), .C(_2266_), );
  OAI21X1 OAI21X1_795 (.Y(_2267_), .A(_2264__bF_buf8), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf4), .C(regs_3__1_), );
  OAI21X1 OAI21X1_796 (.Y(_779_), .A(_2265__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1003__bF_buf0), .C(_2267_), );
  OAI21X1 OAI21X1_797 (.Y(_2268_), .A(_2264__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf3), .C(regs_3__2_), );
  OAI21X1 OAI21X1_798 (.Y(_790_), .A(_2265__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1005__bF_buf0), .C(_2268_), );
  OAI21X1 OAI21X1_799 (.Y(_2269_), .A(_2264__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf2), .C(regs_3__3_), );
  OAI21X1 OAI21X1_800 (.Y(_793_), .A(_2265__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1007__bF_buf0), .C(_2269_), );
  OAI21X1 OAI21X1_801 (.Y(_2270_), .A(_2264__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf1), .C(regs_3__4_), );
  OAI21X1 OAI21X1_802 (.Y(_794_), .A(_2265__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1009__bF_buf3), .C(_2270_), );
  OAI21X1 OAI21X1_803 (.Y(_2271_), .A(_2264__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf0), .C(regs_3__5_), );
  OAI21X1 OAI21X1_804 (.Y(_795_), .A(_2265__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1011__bF_buf3), .C(_2271_), );
  OAI21X1 OAI21X1_805 (.Y(_2272_), .A(_2264__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf5), .C(regs_3__6_), );
  OAI21X1 OAI21X1_806 (.Y(_796_), .A(_2265__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1013__bF_buf3), .C(_2272_), );
  OAI21X1 OAI21X1_807 (.Y(_2273_), .A(_2264__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf4), .C(regs_3__7_), );
  OAI21X1 OAI21X1_808 (.Y(_797_), .A(_2265__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1015__bF_buf3), .C(_2273_), );
  OAI21X1 OAI21X1_809 (.Y(_2274_), .A(_2264__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf3), .C(regs_3__8_), );
  OAI21X1 OAI21X1_810 (.Y(_798_), .A(_2265__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1017__bF_buf3), .C(_2274_), );
  OAI21X1 OAI21X1_811 (.Y(_2275_), .A(_2264__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf2), .C(regs_3__9_), );
  OAI21X1 OAI21X1_812 (.Y(_799_), .A(_2265__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1019__bF_buf3), .C(_2275_), );
  OAI21X1 OAI21X1_813 (.Y(_2276_), .A(_2264__bF_buf10), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf1), .C(regs_3__10_), );
  OAI21X1 OAI21X1_814 (.Y(_769_), .A(_2265__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1021__bF_buf3), .C(_2276_), );
  OAI21X1 OAI21X1_815 (.Y(_2277_), .A(_2264__bF_buf9), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf0), .C(regs_3__11_), );
  OAI21X1 OAI21X1_816 (.Y(_770_), .A(_2265__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1023__bF_buf3), .C(_2277_), );
  OAI21X1 OAI21X1_817 (.Y(_2278_), .A(_2264__bF_buf8), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf5), .C(regs_3__12_), );
  OAI21X1 OAI21X1_818 (.Y(_771_), .A(_2265__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1025__bF_buf3), .C(_2278_), );
  OAI21X1 OAI21X1_819 (.Y(_2279_), .A(_2264__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf4), .C(regs_3__13_), );
  OAI21X1 OAI21X1_820 (.Y(_772_), .A(_2265__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1027__bF_buf3), .C(_2279_), );
  OAI21X1 OAI21X1_821 (.Y(_2280_), .A(_2264__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf3), .C(regs_3__14_), );
  OAI21X1 OAI21X1_822 (.Y(_773_), .A(_2265__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1029__bF_buf3), .C(_2280_), );
  OAI21X1 OAI21X1_823 (.Y(_2281_), .A(_2264__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf2), .C(regs_3__15_), );
  OAI21X1 OAI21X1_824 (.Y(_774_), .A(_2265__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1031__bF_buf3), .C(_2281_), );
  OAI21X1 OAI21X1_825 (.Y(_2282_), .A(_2264__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf1), .C(regs_3__16_), );
  OAI21X1 OAI21X1_826 (.Y(_775_), .A(_2265__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1033__bF_buf3), .C(_2282_), );
  OAI21X1 OAI21X1_827 (.Y(_2283_), .A(_2264__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf0), .C(regs_3__17_), );
  OAI21X1 OAI21X1_828 (.Y(_776_), .A(_2265__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1035__bF_buf3), .C(_2283_), );
  OAI21X1 OAI21X1_829 (.Y(_2284_), .A(_2264__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf5), .C(regs_3__18_), );
  OAI21X1 OAI21X1_830 (.Y(_777_), .A(_2265__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1037__bF_buf3), .C(_2284_), );
  OAI21X1 OAI21X1_831 (.Y(_2285_), .A(_2264__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf4), .C(regs_3__19_), );
  OAI21X1 OAI21X1_832 (.Y(_778_), .A(_2265__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1039__bF_buf3), .C(_2285_), );
  OAI21X1 OAI21X1_833 (.Y(_2286_), .A(_2264__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf3), .C(regs_3__20_), );
  OAI21X1 OAI21X1_834 (.Y(_780_), .A(_2265__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1041__bF_buf3), .C(_2286_), );
  OAI21X1 OAI21X1_835 (.Y(_2287_), .A(_2264__bF_buf10), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf2), .C(regs_3__21_), );
  OAI21X1 OAI21X1_836 (.Y(_781_), .A(_2265__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1043__bF_buf3), .C(_2287_), );
  OAI21X1 OAI21X1_837 (.Y(_2288_), .A(_2264__bF_buf9), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf1), .C(regs_3__22_), );
  OAI21X1 OAI21X1_838 (.Y(_782_), .A(_2265__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1045__bF_buf3), .C(_2288_), );
  OAI21X1 OAI21X1_839 (.Y(_2289_), .A(_2264__bF_buf8), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf0), .C(regs_3__23_), );
  OAI21X1 OAI21X1_840 (.Y(_783_), .A(_2265__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1047__bF_buf3), .C(_2289_), );
  OAI21X1 OAI21X1_841 (.Y(_2290_), .A(_2264__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf5), .C(regs_3__24_), );
  OAI21X1 OAI21X1_842 (.Y(_784_), .A(_2265__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1049__bF_buf3), .C(_2290_), );
  OAI21X1 OAI21X1_843 (.Y(_2291_), .A(_2264__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf4), .C(regs_3__25_), );
  OAI21X1 OAI21X1_844 (.Y(_785_), .A(_2265__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1051__bF_buf3), .C(_2291_), );
  OAI21X1 OAI21X1_845 (.Y(_2292_), .A(_2264__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf3), .C(regs_3__26_), );
  OAI21X1 OAI21X1_846 (.Y(_786_), .A(_2265__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1053__bF_buf3), .C(_2292_), );
  OAI21X1 OAI21X1_847 (.Y(_2293_), .A(_2264__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf2), .C(regs_3__27_), );
  OAI21X1 OAI21X1_848 (.Y(_787_), .A(_2265__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1055__bF_buf3), .C(_2293_), );
  OAI21X1 OAI21X1_849 (.Y(_2294_), .A(_2264__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf1), .C(regs_3__28_), );
  OAI21X1 OAI21X1_850 (.Y(_788_), .A(_2265__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1057__bF_buf3), .C(_2294_), );
  OAI21X1 OAI21X1_851 (.Y(_2295_), .A(_2264__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf0), .C(regs_3__29_), );
  OAI21X1 OAI21X1_852 (.Y(_789_), .A(_2265__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1059__bF_buf3), .C(_2295_), );
  OAI21X1 OAI21X1_853 (.Y(_2296_), .A(_2264__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf5), .C(regs_3__30_), );
  OAI21X1 OAI21X1_854 (.Y(_791_), .A(_2265__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1061__bF_buf3), .C(_2296_), );
  OAI21X1 OAI21X1_855 (.Y(_2297_), .A(_2264__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1142__bF_buf4), .C(regs_3__31_), );
  OAI21X1 OAI21X1_856 (.Y(_792_), .A(_2265__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1063__bF_buf3), .C(_2297_), );
  INVX1 INVX1_1 (.Y(_2298_), .A(_2264__bF_buf10), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_295 (.Y(_2299_), .A(_998_), .gnd(gnd), .vdd(vdd), .B(_2298_), );
  OAI21X1 OAI21X1_857 (.Y(_2300_), .A(_1001__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf9), .C(regs_2__0_), );
  OAI21X1 OAI21X1_858 (.Y(_704_), .A(_2299__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_992__bF_buf3), .C(_2300_), );
  OAI21X1 OAI21X1_859 (.Y(_2301_), .A(_1001__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf8), .C(regs_2__1_), );
  OAI21X1 OAI21X1_860 (.Y(_715_), .A(_2299__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1003__bF_buf3), .C(_2301_), );
  OAI21X1 OAI21X1_861 (.Y(_2302_), .A(_1001__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf7), .C(regs_2__2_), );
  OAI21X1 OAI21X1_862 (.Y(_726_), .A(_2299__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1005__bF_buf3), .C(_2302_), );
  OAI21X1 OAI21X1_863 (.Y(_2303_), .A(_1001__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf6), .C(regs_2__3_), );
  OAI21X1 OAI21X1_864 (.Y(_729_), .A(_2299__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1007__bF_buf3), .C(_2303_), );
  OAI21X1 OAI21X1_865 (.Y(_2304_), .A(_1001__bF_buf9), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf5), .C(regs_2__4_), );
  OAI21X1 OAI21X1_866 (.Y(_730_), .A(_2299__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1009__bF_buf2), .C(_2304_), );
  OAI21X1 OAI21X1_867 (.Y(_2305_), .A(_1001__bF_buf8), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf4), .C(regs_2__5_), );
  OAI21X1 OAI21X1_868 (.Y(_731_), .A(_2299__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1011__bF_buf2), .C(_2305_), );
  OAI21X1 OAI21X1_869 (.Y(_2306_), .A(_1001__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf3), .C(regs_2__6_), );
  OAI21X1 OAI21X1_870 (.Y(_732_), .A(_2299__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1013__bF_buf2), .C(_2306_), );
  OAI21X1 OAI21X1_871 (.Y(_2307_), .A(_1001__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf2), .C(regs_2__7_), );
  OAI21X1 OAI21X1_872 (.Y(_733_), .A(_2299__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1015__bF_buf2), .C(_2307_), );
  OAI21X1 OAI21X1_873 (.Y(_2308_), .A(_1001__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf1), .C(regs_2__8_), );
  OAI21X1 OAI21X1_874 (.Y(_734_), .A(_2299__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1017__bF_buf2), .C(_2308_), );
  OAI21X1 OAI21X1_875 (.Y(_2309_), .A(_1001__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf0), .C(regs_2__9_), );
  OAI21X1 OAI21X1_876 (.Y(_735_), .A(_2299__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1019__bF_buf2), .C(_2309_), );
  OAI21X1 OAI21X1_877 (.Y(_2310_), .A(_1001__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf10), .C(regs_2__10_), );
  OAI21X1 OAI21X1_878 (.Y(_705_), .A(_2299__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1021__bF_buf2), .C(_2310_), );
  OAI21X1 OAI21X1_879 (.Y(_2311_), .A(_1001__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf9), .C(regs_2__11_), );
  OAI21X1 OAI21X1_880 (.Y(_706_), .A(_2299__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1023__bF_buf2), .C(_2311_), );
  OAI21X1 OAI21X1_881 (.Y(_2312_), .A(_1001__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf8), .C(regs_2__12_), );
  OAI21X1 OAI21X1_882 (.Y(_707_), .A(_2299__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1025__bF_buf2), .C(_2312_), );
  OAI21X1 OAI21X1_883 (.Y(_2313_), .A(_1001__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf7), .C(regs_2__13_), );
  OAI21X1 OAI21X1_884 (.Y(_708_), .A(_2299__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1027__bF_buf2), .C(_2313_), );
  OAI21X1 OAI21X1_885 (.Y(_2314_), .A(_1001__bF_buf9), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf6), .C(regs_2__14_), );
  OAI21X1 OAI21X1_886 (.Y(_709_), .A(_2299__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1029__bF_buf2), .C(_2314_), );
  OAI21X1 OAI21X1_887 (.Y(_2315_), .A(_1001__bF_buf8), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf5), .C(regs_2__15_), );
  OAI21X1 OAI21X1_888 (.Y(_710_), .A(_2299__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1031__bF_buf2), .C(_2315_), );
  OAI21X1 OAI21X1_889 (.Y(_2316_), .A(_1001__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf4), .C(regs_2__16_), );
  OAI21X1 OAI21X1_890 (.Y(_711_), .A(_2299__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1033__bF_buf2), .C(_2316_), );
  OAI21X1 OAI21X1_891 (.Y(_2317_), .A(_1001__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf3), .C(regs_2__17_), );
  OAI21X1 OAI21X1_892 (.Y(_712_), .A(_2299__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1035__bF_buf2), .C(_2317_), );
  OAI21X1 OAI21X1_893 (.Y(_2318_), .A(_1001__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf2), .C(regs_2__18_), );
  OAI21X1 OAI21X1_894 (.Y(_713_), .A(_2299__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1037__bF_buf2), .C(_2318_), );
  OAI21X1 OAI21X1_895 (.Y(_2319_), .A(_1001__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf1), .C(regs_2__19_), );
  OAI21X1 OAI21X1_896 (.Y(_714_), .A(_2299__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1039__bF_buf2), .C(_2319_), );
  OAI21X1 OAI21X1_897 (.Y(_2320_), .A(_1001__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf0), .C(regs_2__20_), );
  OAI21X1 OAI21X1_898 (.Y(_716_), .A(_2299__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1041__bF_buf2), .C(_2320_), );
  OAI21X1 OAI21X1_899 (.Y(_2321_), .A(_1001__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf10), .C(regs_2__21_), );
  OAI21X1 OAI21X1_900 (.Y(_717_), .A(_2299__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1043__bF_buf2), .C(_2321_), );
  OAI21X1 OAI21X1_901 (.Y(_2322_), .A(_1001__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf9), .C(regs_2__22_), );
  OAI21X1 OAI21X1_902 (.Y(_718_), .A(_2299__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1045__bF_buf2), .C(_2322_), );
  OAI21X1 OAI21X1_903 (.Y(_2323_), .A(_1001__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf8), .C(regs_2__23_), );
  OAI21X1 OAI21X1_904 (.Y(_719_), .A(_2299__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1047__bF_buf2), .C(_2323_), );
  OAI21X1 OAI21X1_905 (.Y(_2324_), .A(_1001__bF_buf9), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf7), .C(regs_2__24_), );
  OAI21X1 OAI21X1_906 (.Y(_720_), .A(_2299__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1049__bF_buf2), .C(_2324_), );
  OAI21X1 OAI21X1_907 (.Y(_2325_), .A(_1001__bF_buf8), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf6), .C(regs_2__25_), );
  OAI21X1 OAI21X1_908 (.Y(_721_), .A(_2299__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1051__bF_buf2), .C(_2325_), );
  OAI21X1 OAI21X1_909 (.Y(_2326_), .A(_1001__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf5), .C(regs_2__26_), );
  OAI21X1 OAI21X1_910 (.Y(_722_), .A(_2299__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1053__bF_buf2), .C(_2326_), );
  OAI21X1 OAI21X1_911 (.Y(_2327_), .A(_1001__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf4), .C(regs_2__27_), );
  OAI21X1 OAI21X1_912 (.Y(_723_), .A(_2299__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1055__bF_buf2), .C(_2327_), );
  OAI21X1 OAI21X1_913 (.Y(_2328_), .A(_1001__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf3), .C(regs_2__28_), );
  OAI21X1 OAI21X1_914 (.Y(_724_), .A(_2299__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1057__bF_buf2), .C(_2328_), );
  OAI21X1 OAI21X1_915 (.Y(_2329_), .A(_1001__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf2), .C(regs_2__29_), );
  OAI21X1 OAI21X1_916 (.Y(_725_), .A(_2299__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1059__bF_buf2), .C(_2329_), );
  OAI21X1 OAI21X1_917 (.Y(_2330_), .A(_1001__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf1), .C(regs_2__30_), );
  OAI21X1 OAI21X1_918 (.Y(_727_), .A(_2299__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1061__bF_buf2), .C(_2330_), );
  OAI21X1 OAI21X1_919 (.Y(_2331_), .A(_1001__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf0), .C(regs_2__31_), );
  OAI21X1 OAI21X1_920 (.Y(_728_), .A(_2299__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1063__bF_buf2), .C(_2331_), );
  NAND2X1 NAND2X1_296 (.Y(_2332_), .A(_1068_), .gnd(gnd), .vdd(vdd), .B(_2298_), );
  OAI21X1 OAI21X1_921 (.Y(_2333_), .A(_1070__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf10), .C(regs_1__0_), );
  OAI21X1 OAI21X1_922 (.Y(_352_), .A(_2332__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_992__bF_buf2), .C(_2333_), );
  OAI21X1 OAI21X1_923 (.Y(_2334_), .A(_1070__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf9), .C(regs_1__1_), );
  OAI21X1 OAI21X1_924 (.Y(_363_), .A(_2332__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1003__bF_buf2), .C(_2334_), );
  OAI21X1 OAI21X1_925 (.Y(_2335_), .A(_1070__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf8), .C(regs_1__2_), );
  OAI21X1 OAI21X1_926 (.Y(_374_), .A(_2332__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1005__bF_buf2), .C(_2335_), );
  OAI21X1 OAI21X1_927 (.Y(_2336_), .A(_1070__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf7), .C(regs_1__3_), );
  OAI21X1 OAI21X1_928 (.Y(_377_), .A(_2332__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1007__bF_buf2), .C(_2336_), );
  OAI21X1 OAI21X1_929 (.Y(_2337_), .A(_1070__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf6), .C(regs_1__4_), );
  OAI21X1 OAI21X1_930 (.Y(_378_), .A(_2332__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1009__bF_buf1), .C(_2337_), );
  OAI21X1 OAI21X1_931 (.Y(_2338_), .A(_1070__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf5), .C(regs_1__5_), );
  OAI21X1 OAI21X1_932 (.Y(_379_), .A(_2332__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1011__bF_buf1), .C(_2338_), );
  OAI21X1 OAI21X1_933 (.Y(_2339_), .A(_1070__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf4), .C(regs_1__6_), );
  OAI21X1 OAI21X1_934 (.Y(_380_), .A(_2332__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1013__bF_buf1), .C(_2339_), );
  OAI21X1 OAI21X1_935 (.Y(_2340_), .A(_1070__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf3), .C(regs_1__7_), );
  OAI21X1 OAI21X1_936 (.Y(_381_), .A(_2332__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1015__bF_buf1), .C(_2340_), );
  OAI21X1 OAI21X1_937 (.Y(_2341_), .A(_1070__bF_buf10), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf2), .C(regs_1__8_), );
  OAI21X1 OAI21X1_938 (.Y(_382_), .A(_2332__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1017__bF_buf1), .C(_2341_), );
  OAI21X1 OAI21X1_939 (.Y(_2342_), .A(_1070__bF_buf9), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf1), .C(regs_1__9_), );
  OAI21X1 OAI21X1_940 (.Y(_383_), .A(_2332__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1019__bF_buf1), .C(_2342_), );
  OAI21X1 OAI21X1_941 (.Y(_2343_), .A(_1070__bF_buf8), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf0), .C(regs_1__10_), );
  OAI21X1 OAI21X1_942 (.Y(_353_), .A(_2332__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1021__bF_buf1), .C(_2343_), );
  OAI21X1 OAI21X1_943 (.Y(_2344_), .A(_1070__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf10), .C(regs_1__11_), );
  OAI21X1 OAI21X1_944 (.Y(_354_), .A(_2332__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1023__bF_buf1), .C(_2344_), );
  OAI21X1 OAI21X1_945 (.Y(_2345_), .A(_1070__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf9), .C(regs_1__12_), );
  OAI21X1 OAI21X1_946 (.Y(_355_), .A(_2332__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1025__bF_buf1), .C(_2345_), );
  OAI21X1 OAI21X1_947 (.Y(_2346_), .A(_1070__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf8), .C(regs_1__13_), );
  OAI21X1 OAI21X1_948 (.Y(_356_), .A(_2332__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1027__bF_buf1), .C(_2346_), );
  OAI21X1 OAI21X1_949 (.Y(_2347_), .A(_1070__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf7), .C(regs_1__14_), );
  OAI21X1 OAI21X1_950 (.Y(_357_), .A(_2332__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1029__bF_buf1), .C(_2347_), );
  OAI21X1 OAI21X1_951 (.Y(_2348_), .A(_1070__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf6), .C(regs_1__15_), );
  OAI21X1 OAI21X1_952 (.Y(_358_), .A(_2332__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1031__bF_buf1), .C(_2348_), );
  OAI21X1 OAI21X1_953 (.Y(_2349_), .A(_1070__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf5), .C(regs_1__16_), );
  OAI21X1 OAI21X1_954 (.Y(_359_), .A(_2332__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1033__bF_buf1), .C(_2349_), );
  OAI21X1 OAI21X1_955 (.Y(_2350_), .A(_1070__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf4), .C(regs_1__17_), );
  OAI21X1 OAI21X1_956 (.Y(_360_), .A(_2332__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1035__bF_buf1), .C(_2350_), );
  OAI21X1 OAI21X1_957 (.Y(_2351_), .A(_1070__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf3), .C(regs_1__18_), );
  OAI21X1 OAI21X1_958 (.Y(_361_), .A(_2332__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1037__bF_buf1), .C(_2351_), );
  OAI21X1 OAI21X1_959 (.Y(_2352_), .A(_1070__bF_buf10), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf2), .C(regs_1__19_), );
  OAI21X1 OAI21X1_960 (.Y(_362_), .A(_2332__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1039__bF_buf1), .C(_2352_), );
  OAI21X1 OAI21X1_961 (.Y(_2353_), .A(_1070__bF_buf9), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf1), .C(regs_1__20_), );
  OAI21X1 OAI21X1_962 (.Y(_364_), .A(_2332__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1041__bF_buf1), .C(_2353_), );
  OAI21X1 OAI21X1_963 (.Y(_2354_), .A(_1070__bF_buf8), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf0), .C(regs_1__21_), );
  OAI21X1 OAI21X1_964 (.Y(_365_), .A(_2332__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1043__bF_buf1), .C(_2354_), );
  OAI21X1 OAI21X1_965 (.Y(_2355_), .A(_1070__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf10), .C(regs_1__22_), );
  OAI21X1 OAI21X1_966 (.Y(_366_), .A(_2332__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1045__bF_buf1), .C(_2355_), );
  OAI21X1 OAI21X1_967 (.Y(_2356_), .A(_1070__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf9), .C(regs_1__23_), );
  OAI21X1 OAI21X1_968 (.Y(_367_), .A(_2332__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1047__bF_buf1), .C(_2356_), );
  OAI21X1 OAI21X1_969 (.Y(_2357_), .A(_1070__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf8), .C(regs_1__24_), );
  OAI21X1 OAI21X1_970 (.Y(_368_), .A(_2332__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1049__bF_buf1), .C(_2357_), );
  OAI21X1 OAI21X1_971 (.Y(_2358_), .A(_1070__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf7), .C(regs_1__25_), );
  OAI21X1 OAI21X1_972 (.Y(_369_), .A(_2332__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1051__bF_buf1), .C(_2358_), );
  OAI21X1 OAI21X1_973 (.Y(_2359_), .A(_1070__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf6), .C(regs_1__26_), );
  OAI21X1 OAI21X1_974 (.Y(_370_), .A(_2332__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1053__bF_buf1), .C(_2359_), );
  OAI21X1 OAI21X1_975 (.Y(_2360_), .A(_1070__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf5), .C(regs_1__27_), );
  OAI21X1 OAI21X1_976 (.Y(_371_), .A(_2332__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1055__bF_buf1), .C(_2360_), );
  OAI21X1 OAI21X1_977 (.Y(_2361_), .A(_1070__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf4), .C(regs_1__28_), );
  OAI21X1 OAI21X1_978 (.Y(_372_), .A(_2332__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1057__bF_buf1), .C(_2361_), );
  OAI21X1 OAI21X1_979 (.Y(_2362_), .A(_1070__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf3), .C(regs_1__29_), );
  OAI21X1 OAI21X1_980 (.Y(_373_), .A(_2332__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1059__bF_buf1), .C(_2362_), );
  OAI21X1 OAI21X1_981 (.Y(_2363_), .A(_1070__bF_buf10), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf2), .C(regs_1__30_), );
  OAI21X1 OAI21X1_982 (.Y(_375_), .A(_2332__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1061__bF_buf1), .C(_2363_), );
  OAI21X1 OAI21X1_983 (.Y(_2364_), .A(_1070__bF_buf9), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf1), .C(regs_1__31_), );
  OAI21X1 OAI21X1_984 (.Y(_376_), .A(_2332__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1063__bF_buf1), .C(_2364_), );
  NAND2X1 NAND2X1_297 (.Y(_2365_), .A(_1273_), .gnd(gnd), .vdd(vdd), .B(_2298_), );
  OAI21X1 OAI21X1_985 (.Y(_2366_), .A(_1104__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf0), .C(regs_0__0_), );
  OAI21X1 OAI21X1_986 (.Y(_0_), .A(_2365__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_992__bF_buf1), .C(_2366_), );
  OAI21X1 OAI21X1_987 (.Y(_2367_), .A(_1104__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf10), .C(regs_0__1_), );
  OAI21X1 OAI21X1_988 (.Y(_11_), .A(_2365__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1003__bF_buf1), .C(_2367_), );
  OAI21X1 OAI21X1_989 (.Y(_2368_), .A(_1104__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf9), .C(regs_0__2_), );
  OAI21X1 OAI21X1_990 (.Y(_22_), .A(_2365__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1005__bF_buf1), .C(_2368_), );
  OAI21X1 OAI21X1_991 (.Y(_2369_), .A(_1104__bF_buf14), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf8), .C(regs_0__3_), );
  OAI21X1 OAI21X1_992 (.Y(_25_), .A(_2365__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1007__bF_buf1), .C(_2369_), );
  OAI21X1 OAI21X1_993 (.Y(_2370_), .A(_1104__bF_buf13), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf7), .C(regs_0__4_), );
  OAI21X1 OAI21X1_994 (.Y(_26_), .A(_2365__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1009__bF_buf0), .C(_2370_), );
  OAI21X1 OAI21X1_995 (.Y(_2371_), .A(_1104__bF_buf12), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf6), .C(regs_0__5_), );
  OAI21X1 OAI21X1_996 (.Y(_27_), .A(_2365__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1011__bF_buf0), .C(_2371_), );
  OAI21X1 OAI21X1_997 (.Y(_2372_), .A(_1104__bF_buf11), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf5), .C(regs_0__6_), );
  OAI21X1 OAI21X1_998 (.Y(_28_), .A(_2365__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1013__bF_buf0), .C(_2372_), );
  OAI21X1 OAI21X1_999 (.Y(_2373_), .A(_1104__bF_buf10), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf4), .C(regs_0__7_), );
  OAI21X1 OAI21X1_1000 (.Y(_29_), .A(_2365__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1015__bF_buf0), .C(_2373_), );
  OAI21X1 OAI21X1_1001 (.Y(_2374_), .A(_1104__bF_buf9), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf3), .C(regs_0__8_), );
  OAI21X1 OAI21X1_1002 (.Y(_30_), .A(_2365__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1017__bF_buf0), .C(_2374_), );
  OAI21X1 OAI21X1_1003 (.Y(_2375_), .A(_1104__bF_buf8), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf2), .C(regs_0__9_), );
  OAI21X1 OAI21X1_1004 (.Y(_31_), .A(_2365__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1019__bF_buf0), .C(_2375_), );
  OAI21X1 OAI21X1_1005 (.Y(_2376_), .A(_1104__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf1), .C(regs_0__10_), );
  OAI21X1 OAI21X1_1006 (.Y(_1_), .A(_2365__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1021__bF_buf0), .C(_2376_), );
  OAI21X1 OAI21X1_1007 (.Y(_2377_), .A(_1104__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf0), .C(regs_0__11_), );
  OAI21X1 OAI21X1_1008 (.Y(_2_), .A(_2365__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1023__bF_buf0), .C(_2377_), );
  OAI21X1 OAI21X1_1009 (.Y(_2378_), .A(_1104__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf10), .C(regs_0__12_), );
  OAI21X1 OAI21X1_1010 (.Y(_3_), .A(_2365__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1025__bF_buf0), .C(_2378_), );
  OAI21X1 OAI21X1_1011 (.Y(_2379_), .A(_1104__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf9), .C(regs_0__13_), );
  OAI21X1 OAI21X1_1012 (.Y(_4_), .A(_2365__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1027__bF_buf0), .C(_2379_), );
  OAI21X1 OAI21X1_1013 (.Y(_2380_), .A(_1104__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf8), .C(regs_0__14_), );
  OAI21X1 OAI21X1_1014 (.Y(_5_), .A(_2365__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1029__bF_buf0), .C(_2380_), );
  OAI21X1 OAI21X1_1015 (.Y(_2381_), .A(_1104__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf7), .C(regs_0__15_), );
  OAI21X1 OAI21X1_1016 (.Y(_6_), .A(_2365__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1031__bF_buf0), .C(_2381_), );
  OAI21X1 OAI21X1_1017 (.Y(_2382_), .A(_1104__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf6), .C(regs_0__16_), );
  OAI21X1 OAI21X1_1018 (.Y(_7_), .A(_2365__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1033__bF_buf0), .C(_2382_), );
  OAI21X1 OAI21X1_1019 (.Y(_2383_), .A(_1104__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf5), .C(regs_0__17_), );
  OAI21X1 OAI21X1_1020 (.Y(_8_), .A(_2365__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1035__bF_buf0), .C(_2383_), );
  OAI21X1 OAI21X1_1021 (.Y(_2384_), .A(_1104__bF_buf14), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf4), .C(regs_0__18_), );
  OAI21X1 OAI21X1_1022 (.Y(_9_), .A(_2365__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1037__bF_buf0), .C(_2384_), );
  OAI21X1 OAI21X1_1023 (.Y(_2385_), .A(_1104__bF_buf13), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf3), .C(regs_0__19_), );
  OAI21X1 OAI21X1_1024 (.Y(_10_), .A(_2365__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1039__bF_buf0), .C(_2385_), );
  OAI21X1 OAI21X1_1025 (.Y(_2386_), .A(_1104__bF_buf12), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf2), .C(regs_0__20_), );
  OAI21X1 OAI21X1_1026 (.Y(_12_), .A(_2365__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1041__bF_buf0), .C(_2386_), );
  OAI21X1 OAI21X1_1027 (.Y(_2387_), .A(_1104__bF_buf11), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf1), .C(regs_0__21_), );
  OAI21X1 OAI21X1_1028 (.Y(_13_), .A(_2365__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1043__bF_buf0), .C(_2387_), );
  OAI21X1 OAI21X1_1029 (.Y(_2388_), .A(_1104__bF_buf10), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf0), .C(regs_0__22_), );
  OAI21X1 OAI21X1_1030 (.Y(_14_), .A(_2365__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1045__bF_buf0), .C(_2388_), );
  OAI21X1 OAI21X1_1031 (.Y(_2389_), .A(_1104__bF_buf9), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf10), .C(regs_0__23_), );
  OAI21X1 OAI21X1_1032 (.Y(_15_), .A(_2365__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1047__bF_buf0), .C(_2389_), );
  OAI21X1 OAI21X1_1033 (.Y(_2390_), .A(_1104__bF_buf8), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf9), .C(regs_0__24_), );
  OAI21X1 OAI21X1_1034 (.Y(_16_), .A(_2365__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1049__bF_buf0), .C(_2390_), );
  OAI21X1 OAI21X1_1035 (.Y(_2391_), .A(_1104__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf8), .C(regs_0__25_), );
  OAI21X1 OAI21X1_1036 (.Y(_17_), .A(_2365__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1051__bF_buf0), .C(_2391_), );
  OAI21X1 OAI21X1_1037 (.Y(_2392_), .A(_1104__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf7), .C(regs_0__26_), );
  OAI21X1 OAI21X1_1038 (.Y(_18_), .A(_2365__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1053__bF_buf0), .C(_2392_), );
  OAI21X1 OAI21X1_1039 (.Y(_2393_), .A(_1104__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf6), .C(regs_0__27_), );
  OAI21X1 OAI21X1_1040 (.Y(_19_), .A(_2365__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_1055__bF_buf0), .C(_2393_), );
  OAI21X1 OAI21X1_1041 (.Y(_2394_), .A(_1104__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf5), .C(regs_0__28_), );
  OAI21X1 OAI21X1_1042 (.Y(_20_), .A(_2365__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_1057__bF_buf0), .C(_2394_), );
  OAI21X1 OAI21X1_1043 (.Y(_2395_), .A(_1104__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf4), .C(regs_0__29_), );
  OAI21X1 OAI21X1_1044 (.Y(_21_), .A(_2365__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_1059__bF_buf0), .C(_2395_), );
  OAI21X1 OAI21X1_1045 (.Y(_2396_), .A(_1104__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf3), .C(regs_0__30_), );
  OAI21X1 OAI21X1_1046 (.Y(_23_), .A(_2365__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_1061__bF_buf0), .C(_2396_), );
  OAI21X1 OAI21X1_1047 (.Y(_2397_), .A(_1104__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_2264__bF_buf2), .C(regs_0__31_), );
  OAI21X1 OAI21X1_1048 (.Y(_24_), .A(_2365__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_1063__bF_buf0), .C(_2397_), );
  INVX8 INVX8_2 (.Y(_2398_), .A(raddr1[3]), .gnd(gnd), .vdd(vdd), );
  INVX8 INVX8_3 (.Y(_2399_), .A(raddr1_2_bF_buf10_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_298 (.Y(_2400_), .A(regs_22__0_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf96_), );
  OAI21X1 OAI21X1_1049 (.Y(_2401_), .A(_1307_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf95_), .C(_2400_), );
  NAND2X1 NAND2X1_299 (.Y(_2402_), .A(regs_20__0_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf94_), );
  OAI21X1 OAI21X1_1050 (.Y(_2403_), .A(_1407_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf93_), .C(_2402_), );
  MUX2X1 MUX2X1_1 (.Y(_2404_), .A(_2403_), .gnd(gnd), .vdd(vdd), .B(_2401_), .S(raddr1_1_bF_buf14_bF_buf3_), );
  NAND2X1 NAND2X1_300 (.Y(_2405_), .A(_2399__bF_buf8), .gnd(gnd), .vdd(vdd), .B(_2404_), );
  NAND2X1 NAND2X1_301 (.Y(_2406_), .A(regs_18__0_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf92_), );
  OAI21X1 OAI21X1_1051 (.Y(_2407_), .A(_1505_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf91_), .C(_2406_), );
  NAND2X1 NAND2X1_302 (.Y(_2408_), .A(regs_16__0_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf90_), );
  OAI21X1 OAI21X1_1052 (.Y(_2409_), .A(_1604_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf89_), .C(_2408_), );
  MUX2X1 MUX2X1_2 (.Y(_2410_), .A(_2409_), .gnd(gnd), .vdd(vdd), .B(_2407_), .S(raddr1_1_bF_buf13_bF_buf3_), );
  AOI21X1 AOI21X1_129 (.Y(_2411_), .A(raddr1_2_bF_buf9_), .gnd(gnd), .vdd(vdd), .B(_2410_), .C(_2398__bF_buf7), );
  AND2X2 AND2X2_1 (.Y(_2412_), .A(regs_26__0_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf88_), );
  OAI21X1 OAI21X1_1053 (.Y(_2413_), .A(_1138_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf87_), .C(raddr1_2_bF_buf8_), );
  NOR2X1 NOR2X1_143 (.Y(_2414_), .A(_2412_), .gnd(gnd), .vdd(vdd), .B(_2413_), );
  INVX8 INVX8_4 (.Y(_2415_), .A(raddr1_1_bF_buf12_bF_buf3_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1054 (.Y(_2416_), .A(regs_30__0_), .gnd(gnd), .vdd(vdd), .B(raddr1_2_bF_buf7_), .C(_2415__bF_buf8), );
  INVX1 INVX1_2 (.Y(_2417_), .A(regs_25__0_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1055 (.Y(_2418_), .A(_2417_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf86_), .C(raddr1_2_bF_buf6_), );
  AOI21X1 AOI21X1_130 (.Y(_2419_), .A(regs_24__0_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf85_), .C(_2418_), );
  INVX1 INVX1_3 (.Y(_2420_), .A(regs_29__0_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_144 (.Y(_2421_), .A(raddr1_0_bF_buf84_), .gnd(gnd), .vdd(vdd), .B(_2420_), );
  NAND2X1 NAND2X1_303 (.Y(_2422_), .A(regs_28__0_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf83_), );
  NAND2X1 NAND2X1_304 (.Y(_2423_), .A(_2399__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_2422_), );
  OAI21X1 OAI21X1_1056 (.Y(_2424_), .A(_2423_), .gnd(gnd), .vdd(vdd), .B(_2421_), .C(raddr1_1_bF_buf11_bF_buf3_), );
  OAI22X1 OAI22X1_1 (.Y(_2425_), .A(_2414_), .gnd(gnd), .vdd(vdd), .B(_2416_), .C(_2424_), .D(_2419_), );
  AOI22X1 AOI22X1_1 (.Y(_2426_), .A(_2425_), .gnd(gnd), .vdd(vdd), .B(_2398__bF_buf6), .C(_2405_), .D(_2411_), );
  INVX1 INVX1_4 (.Y(_2427_), .A(regs_5__0_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1057 (.Y(_2428_), .A(_2427_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf82_), .C(raddr1_1_bF_buf10_bF_buf3_), );
  AOI21X1 AOI21X1_131 (.Y(_2429_), .A(regs_4__0_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf81_), .C(_2428_), );
  AND2X2 AND2X2_2 (.Y(_2430_), .A(regs_6__0_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf80_), );
  OAI21X1 OAI21X1_1058 (.Y(_2431_), .A(_2097_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf79_), .C(_2415__bF_buf7), );
  OAI21X1 OAI21X1_1059 (.Y(_2432_), .A(_2431_), .gnd(gnd), .vdd(vdd), .B(_2430_), .C(_2399__bF_buf6), );
  INVX1 INVX1_5 (.Y(_2433_), .A(regs_1__0_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1060 (.Y(_2434_), .A(_2433_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf78_), .C(raddr1_1_bF_buf9_bF_buf3_), );
  AOI21X1 AOI21X1_132 (.Y(_2435_), .A(regs_0__0_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf77_), .C(_2434_), );
  INVX1 INVX1_6 (.Y(_2436_), .A(regs_3__0_), .gnd(gnd), .vdd(vdd), );
  AOI21X1 AOI21X1_133 (.Y(_2437_), .A(regs_2__0_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf76_), .C(raddr1_1_bF_buf8_), );
  OAI21X1 OAI21X1_1061 (.Y(_2438_), .A(_2436_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf75_), .C(_2437_), );
  NAND2X1 NAND2X1_305 (.Y(_2439_), .A(raddr1_2_bF_buf5_), .gnd(gnd), .vdd(vdd), .B(_2438_), );
  OAI22X1 OAI22X1_2 (.Y(_2440_), .A(_2439_), .gnd(gnd), .vdd(vdd), .B(_2435_), .C(_2432_), .D(_2429_), );
  NAND2X1 NAND2X1_306 (.Y(_2441_), .A(regs_10__0_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf74_), );
  OAI21X1 OAI21X1_1062 (.Y(_2442_), .A(_1900_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf73_), .C(_2441_), );
  NAND2X1 NAND2X1_307 (.Y(_2443_), .A(regs_8__0_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf72_), );
  OAI21X1 OAI21X1_1063 (.Y(_2444_), .A(_1999_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf71_), .C(_2443_), );
  MUX2X1 MUX2X1_3 (.Y(_2445_), .A(_2444_), .gnd(gnd), .vdd(vdd), .B(_2442_), .S(raddr1_1_bF_buf7_), );
  NAND2X1 NAND2X1_308 (.Y(_2446_), .A(regs_14__0_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf70_), );
  OAI21X1 OAI21X1_1064 (.Y(_2447_), .A(_1702_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf69_), .C(_2446_), );
  NAND2X1 NAND2X1_309 (.Y(_2448_), .A(regs_12__0_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf68_), );
  OAI21X1 OAI21X1_1065 (.Y(_2449_), .A(_1802_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf67_), .C(_2448_), );
  MUX2X1 MUX2X1_4 (.Y(_2450_), .A(_2449_), .gnd(gnd), .vdd(vdd), .B(_2447_), .S(raddr1_1_bF_buf6_), );
  MUX2X1 MUX2X1_5 (.Y(_2451_), .A(_2450_), .gnd(gnd), .vdd(vdd), .B(_2445_), .S(_2399__bF_buf5), );
  MUX2X1 MUX2X1_6 (.Y(_2452_), .A(_2451_), .gnd(gnd), .vdd(vdd), .B(_2440_), .S(_2398__bF_buf5), );
  MUX2X1 MUX2X1_7 (.Y(_5511__0_), .A(_2452_), .gnd(gnd), .vdd(vdd), .B(_2426_), .S(raddr1_4_bF_buf4_), );
  OAI21X1 OAI21X1_1066 (.Y(_2453_), .A(_1410_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf66_), .C(raddr1_1_bF_buf5_), );
  AOI21X1 AOI21X1_134 (.Y(_2454_), .A(regs_20__1_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf65_), .C(_2453_), );
  AND2X2 AND2X2_3 (.Y(_2455_), .A(regs_22__1_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf64_), );
  OAI21X1 OAI21X1_1067 (.Y(_2456_), .A(_1312_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf63_), .C(_2415__bF_buf6), );
  OAI21X1 OAI21X1_1068 (.Y(_2457_), .A(_2456_), .gnd(gnd), .vdd(vdd), .B(_2455_), .C(_2399__bF_buf4), );
  OAI21X1 OAI21X1_1069 (.Y(_2458_), .A(_1607_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf62_), .C(raddr1_1_bF_buf4_), );
  AOI21X1 AOI21X1_135 (.Y(_2459_), .A(regs_16__1_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf61_), .C(_2458_), );
  NOR2X1 NOR2X1_145 (.Y(_2460_), .A(raddr1_0_bF_buf60_), .gnd(gnd), .vdd(vdd), .B(_1509_), );
  NAND2X1 NAND2X1_310 (.Y(_2461_), .A(regs_18__1_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf59_), );
  NAND2X1 NAND2X1_311 (.Y(_2462_), .A(_2415__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_2461_), );
  OAI21X1 OAI21X1_1070 (.Y(_2463_), .A(_2462_), .gnd(gnd), .vdd(vdd), .B(_2460_), .C(raddr1_2_bF_buf4_), );
  OAI22X1 OAI22X1_3 (.Y(_2464_), .A(_2459_), .gnd(gnd), .vdd(vdd), .B(_2463_), .C(_2457_), .D(_2454_), );
  INVX1 INVX1_7 (.Y(_2465_), .A(regs_29__1_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_312 (.Y(_2466_), .A(regs_28__1_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf58_), );
  OAI21X1 OAI21X1_1071 (.Y(_2467_), .A(_2465_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf57_), .C(_2466_), );
  MUX2X1 MUX2X1_8 (.Y(_2468_), .A(_2467_), .gnd(gnd), .vdd(vdd), .B(regs_30__1_), .S(raddr1_1_bF_buf3_), );
  NAND2X1 NAND2X1_313 (.Y(_2469_), .A(regs_26__1_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf56_), );
  OAI21X1 OAI21X1_1072 (.Y(_2470_), .A(_1145_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf55_), .C(_2469_), );
  INVX1 INVX1_8 (.Y(_2471_), .A(regs_25__1_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_314 (.Y(_2472_), .A(regs_24__1_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf54_), );
  OAI21X1 OAI21X1_1073 (.Y(_2473_), .A(_2471_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf53_), .C(_2472_), );
  MUX2X1 MUX2X1_9 (.Y(_2474_), .A(_2473_), .gnd(gnd), .vdd(vdd), .B(_2470_), .S(raddr1_1_bF_buf2_), );
  MUX2X1 MUX2X1_10 (.Y(_2475_), .A(_2474_), .gnd(gnd), .vdd(vdd), .B(_2468_), .S(raddr1_2_bF_buf3_), );
  MUX2X1 MUX2X1_11 (.Y(_2476_), .A(_2475_), .gnd(gnd), .vdd(vdd), .B(_2464_), .S(_2398__bF_buf4), );
  NAND2X1 NAND2X1_315 (.Y(_2477_), .A(regs_6__1_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf52_), );
  OAI21X1 OAI21X1_1074 (.Y(_2478_), .A(_2103_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf51_), .C(_2477_), );
  INVX1 INVX1_9 (.Y(_2479_), .A(regs_5__1_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_316 (.Y(_2480_), .A(regs_4__1_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf50_), );
  OAI21X1 OAI21X1_1075 (.Y(_2481_), .A(_2479_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf49_), .C(_2480_), );
  MUX2X1 MUX2X1_12 (.Y(_2482_), .A(_2481_), .gnd(gnd), .vdd(vdd), .B(_2478_), .S(raddr1_1_bF_buf1_), );
  INVX1 INVX1_10 (.Y(_2483_), .A(regs_3__1_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_317 (.Y(_2484_), .A(regs_2__1_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf48_), );
  OAI21X1 OAI21X1_1076 (.Y(_2485_), .A(_2483_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf47_), .C(_2484_), );
  INVX1 INVX1_11 (.Y(_2486_), .A(regs_1__1_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_318 (.Y(_2487_), .A(regs_0__1_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf46_), );
  OAI21X1 OAI21X1_1077 (.Y(_2488_), .A(_2486_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf45_), .C(_2487_), );
  MUX2X1 MUX2X1_13 (.Y(_2489_), .A(_2488_), .gnd(gnd), .vdd(vdd), .B(_2485_), .S(raddr1_1_bF_buf0_), );
  MUX2X1 MUX2X1_14 (.Y(_2490_), .A(_2489_), .gnd(gnd), .vdd(vdd), .B(_2482_), .S(raddr1_2_bF_buf2_), );
  NAND2X1 NAND2X1_319 (.Y(_2491_), .A(regs_10__1_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf44_), );
  OAI21X1 OAI21X1_1078 (.Y(_2492_), .A(_1904_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf43_), .C(_2491_), );
  NAND2X1 NAND2X1_320 (.Y(_2493_), .A(regs_8__1_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf42_), );
  OAI21X1 OAI21X1_1079 (.Y(_2494_), .A(_2002_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf41_), .C(_2493_), );
  MUX2X1 MUX2X1_15 (.Y(_2495_), .A(_2494_), .gnd(gnd), .vdd(vdd), .B(_2492_), .S(raddr1_1_bF_buf14_bF_buf2_), );
  NAND2X1 NAND2X1_321 (.Y(_2496_), .A(regs_14__1_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf40_), );
  OAI21X1 OAI21X1_1080 (.Y(_2497_), .A(_1707_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf39_), .C(_2496_), );
  NAND2X1 NAND2X1_322 (.Y(_2498_), .A(regs_12__1_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf38_), );
  OAI21X1 OAI21X1_1081 (.Y(_2499_), .A(_1805_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf37_), .C(_2498_), );
  MUX2X1 MUX2X1_16 (.Y(_2500_), .A(_2499_), .gnd(gnd), .vdd(vdd), .B(_2497_), .S(raddr1_1_bF_buf13_bF_buf2_), );
  MUX2X1 MUX2X1_17 (.Y(_2501_), .A(_2500_), .gnd(gnd), .vdd(vdd), .B(_2495_), .S(_2399__bF_buf3), );
  MUX2X1 MUX2X1_18 (.Y(_2502_), .A(_2501_), .gnd(gnd), .vdd(vdd), .B(_2490_), .S(_2398__bF_buf3), );
  MUX2X1 MUX2X1_19 (.Y(_5511__1_), .A(_2502_), .gnd(gnd), .vdd(vdd), .B(_2476_), .S(raddr1_4_bF_buf3_), );
  NAND2X1 NAND2X1_323 (.Y(_2503_), .A(regs_22__2_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf36_), );
  OAI21X1 OAI21X1_1082 (.Y(_2504_), .A(_1314_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf35_), .C(_2503_), );
  NAND2X1 NAND2X1_324 (.Y(_2505_), .A(regs_20__2_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf34_), );
  OAI21X1 OAI21X1_1083 (.Y(_2506_), .A(_1412_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf33_), .C(_2505_), );
  MUX2X1 MUX2X1_20 (.Y(_2507_), .A(_2506_), .gnd(gnd), .vdd(vdd), .B(_2504_), .S(raddr1_1_bF_buf12_bF_buf2_), );
  NAND2X1 NAND2X1_325 (.Y(_2508_), .A(_2399__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_2507_), );
  NAND2X1 NAND2X1_326 (.Y(_2509_), .A(regs_18__2_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf32_), );
  OAI21X1 OAI21X1_1084 (.Y(_2510_), .A(_1511_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf31_), .C(_2509_), );
  NAND2X1 NAND2X1_327 (.Y(_2511_), .A(regs_16__2_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf30_), );
  OAI21X1 OAI21X1_1085 (.Y(_2512_), .A(_1609_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf29_), .C(_2511_), );
  MUX2X1 MUX2X1_21 (.Y(_2513_), .A(_2512_), .gnd(gnd), .vdd(vdd), .B(_2510_), .S(raddr1_1_bF_buf11_bF_buf2_), );
  AOI21X1 AOI21X1_136 (.Y(_2514_), .A(raddr1_2_bF_buf1_), .gnd(gnd), .vdd(vdd), .B(_2513_), .C(_2398__bF_buf2), );
  OAI21X1 OAI21X1_1086 (.Y(_2515_), .A(_1147_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf28_), .C(raddr1_2_bF_buf0_), );
  AOI21X1 AOI21X1_137 (.Y(_2516_), .A(regs_26__2_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf27_), .C(_2515_), );
  OAI21X1 OAI21X1_1087 (.Y(_2517_), .A(regs_30__2_), .gnd(gnd), .vdd(vdd), .B(raddr1_2_bF_buf10_), .C(_2415__bF_buf4), );
  INVX1 INVX1_12 (.Y(_2518_), .A(regs_25__2_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1088 (.Y(_2519_), .A(_2518_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf26_), .C(raddr1_2_bF_buf9_), );
  AOI21X1 AOI21X1_138 (.Y(_2520_), .A(regs_24__2_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf25_), .C(_2519_), );
  INVX1 INVX1_13 (.Y(_2521_), .A(regs_29__2_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_146 (.Y(_2522_), .A(raddr1_0_bF_buf24_), .gnd(gnd), .vdd(vdd), .B(_2521_), );
  NAND2X1 NAND2X1_328 (.Y(_2523_), .A(regs_28__2_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf23_), );
  NAND2X1 NAND2X1_329 (.Y(_2524_), .A(_2399__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_2523_), );
  OAI21X1 OAI21X1_1089 (.Y(_2525_), .A(_2524_), .gnd(gnd), .vdd(vdd), .B(_2522_), .C(raddr1_1_bF_buf10_bF_buf2_), );
  OAI22X1 OAI22X1_4 (.Y(_2526_), .A(_2516_), .gnd(gnd), .vdd(vdd), .B(_2517_), .C(_2525_), .D(_2520_), );
  AOI22X1 AOI22X1_2 (.Y(_2527_), .A(_2526_), .gnd(gnd), .vdd(vdd), .B(_2398__bF_buf1), .C(_2508_), .D(_2514_), );
  NAND2X1 NAND2X1_330 (.Y(_2528_), .A(regs_6__2_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf22_), );
  OAI21X1 OAI21X1_1090 (.Y(_2529_), .A(_2105_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf21_), .C(_2528_), );
  INVX1 INVX1_14 (.Y(_2530_), .A(regs_5__2_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_331 (.Y(_2531_), .A(regs_4__2_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf20_), );
  OAI21X1 OAI21X1_1091 (.Y(_2532_), .A(_2530_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf19_), .C(_2531_), );
  MUX2X1 MUX2X1_22 (.Y(_2533_), .A(_2532_), .gnd(gnd), .vdd(vdd), .B(_2529_), .S(raddr1_1_bF_buf9_bF_buf2_), );
  INVX1 INVX1_15 (.Y(_2534_), .A(regs_3__2_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_332 (.Y(_2535_), .A(regs_2__2_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf18_), );
  OAI21X1 OAI21X1_1092 (.Y(_2536_), .A(_2534_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf17_), .C(_2535_), );
  INVX1 INVX1_16 (.Y(_2537_), .A(regs_1__2_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_333 (.Y(_2538_), .A(regs_0__2_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf16_), );
  OAI21X1 OAI21X1_1093 (.Y(_2539_), .A(_2537_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf15_), .C(_2538_), );
  MUX2X1 MUX2X1_23 (.Y(_2540_), .A(_2539_), .gnd(gnd), .vdd(vdd), .B(_2536_), .S(raddr1_1_bF_buf8_), );
  MUX2X1 MUX2X1_24 (.Y(_2541_), .A(_2540_), .gnd(gnd), .vdd(vdd), .B(_2533_), .S(raddr1_2_bF_buf8_), );
  NAND2X1 NAND2X1_334 (.Y(_2542_), .A(regs_14__2_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf14_), );
  OAI21X1 OAI21X1_1094 (.Y(_2543_), .A(_1709_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf13_), .C(_2542_), );
  NAND2X1 NAND2X1_335 (.Y(_2544_), .A(regs_12__2_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf12_), );
  OAI21X1 OAI21X1_1095 (.Y(_2545_), .A(_1807_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf11_), .C(_2544_), );
  MUX2X1 MUX2X1_25 (.Y(_2546_), .A(_2545_), .gnd(gnd), .vdd(vdd), .B(_2543_), .S(raddr1_1_bF_buf7_), );
  NAND2X1 NAND2X1_336 (.Y(_2547_), .A(regs_10__2_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf10_), );
  OAI21X1 OAI21X1_1096 (.Y(_2548_), .A(_1906_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf9_), .C(_2547_), );
  NAND2X1 NAND2X1_337 (.Y(_2549_), .A(regs_8__2_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf8_), );
  OAI21X1 OAI21X1_1097 (.Y(_2550_), .A(_2004_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf7_), .C(_2549_), );
  MUX2X1 MUX2X1_26 (.Y(_2551_), .A(_2550_), .gnd(gnd), .vdd(vdd), .B(_2548_), .S(raddr1_1_bF_buf6_), );
  MUX2X1 MUX2X1_27 (.Y(_2552_), .A(_2551_), .gnd(gnd), .vdd(vdd), .B(_2546_), .S(raddr1_2_bF_buf7_), );
  MUX2X1 MUX2X1_28 (.Y(_2553_), .A(_2552_), .gnd(gnd), .vdd(vdd), .B(_2541_), .S(_2398__bF_buf0), );
  MUX2X1 MUX2X1_29 (.Y(_5511__2_), .A(_2553_), .gnd(gnd), .vdd(vdd), .B(_2527_), .S(raddr1_4_bF_buf2_), );
  INVX1 INVX1_17 (.Y(_2554_), .A(regs_5__3_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1098 (.Y(_2555_), .A(_2554_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf6_), .C(raddr1_1_bF_buf5_), );
  AOI21X1 AOI21X1_139 (.Y(_2556_), .A(regs_4__3_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf5_), .C(_2555_), );
  AND2X2 AND2X2_4 (.Y(_2557_), .A(regs_6__3_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf4_), );
  OAI21X1 OAI21X1_1099 (.Y(_2558_), .A(_2107_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf3_), .C(_2415__bF_buf3), );
  OAI21X1 OAI21X1_1100 (.Y(_2559_), .A(_2558_), .gnd(gnd), .vdd(vdd), .B(_2557_), .C(_2399__bF_buf0), );
  INVX1 INVX1_18 (.Y(_2560_), .A(regs_1__3_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1101 (.Y(_2561_), .A(_2560_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf2_), .C(raddr1_1_bF_buf4_), );
  AOI21X1 AOI21X1_140 (.Y(_2562_), .A(regs_0__3_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf1_), .C(_2561_), );
  INVX1 INVX1_19 (.Y(_2563_), .A(regs_3__3_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_147 (.Y(_2564_), .A(raddr1_0_bF_buf0_), .gnd(gnd), .vdd(vdd), .B(_2563_), );
  NAND2X1 NAND2X1_338 (.Y(_2565_), .A(regs_2__3_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf96_), );
  NAND2X1 NAND2X1_339 (.Y(_2566_), .A(_2415__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_2565_), );
  OAI21X1 OAI21X1_1102 (.Y(_2567_), .A(_2566_), .gnd(gnd), .vdd(vdd), .B(_2564_), .C(raddr1_2_bF_buf6_), );
  OAI22X1 OAI22X1_5 (.Y(_2568_), .A(_2562_), .gnd(gnd), .vdd(vdd), .B(_2567_), .C(_2559_), .D(_2556_), );
  NAND2X1 NAND2X1_340 (.Y(_2569_), .A(regs_10__3_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf95_), );
  OAI21X1 OAI21X1_1103 (.Y(_2570_), .A(_1908_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf94_), .C(_2569_), );
  NAND2X1 NAND2X1_341 (.Y(_2571_), .A(regs_8__3_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf93_), );
  OAI21X1 OAI21X1_1104 (.Y(_2572_), .A(_2006_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf92_), .C(_2571_), );
  MUX2X1 MUX2X1_30 (.Y(_2573_), .A(_2572_), .gnd(gnd), .vdd(vdd), .B(_2570_), .S(raddr1_1_bF_buf3_), );
  NAND2X1 NAND2X1_342 (.Y(_2574_), .A(regs_14__3_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf91_), );
  OAI21X1 OAI21X1_1105 (.Y(_2575_), .A(_1711_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf90_), .C(_2574_), );
  NAND2X1 NAND2X1_343 (.Y(_2576_), .A(regs_12__3_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf89_), );
  OAI21X1 OAI21X1_1106 (.Y(_2577_), .A(_1809_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf88_), .C(_2576_), );
  MUX2X1 MUX2X1_31 (.Y(_2578_), .A(_2577_), .gnd(gnd), .vdd(vdd), .B(_2575_), .S(raddr1_1_bF_buf2_), );
  MUX2X1 MUX2X1_32 (.Y(_2579_), .A(_2578_), .gnd(gnd), .vdd(vdd), .B(_2573_), .S(_2399__bF_buf8), );
  MUX2X1 MUX2X1_33 (.Y(_2580_), .A(_2579_), .gnd(gnd), .vdd(vdd), .B(_2568_), .S(_2398__bF_buf7), );
  OAI21X1 OAI21X1_1107 (.Y(_2581_), .A(_1611_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf87_), .C(raddr1_1_bF_buf1_), );
  AOI21X1 AOI21X1_141 (.Y(_2582_), .A(regs_16__3_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf86_), .C(_2581_), );
  NOR2X1 NOR2X1_148 (.Y(_2583_), .A(raddr1_0_bF_buf85_), .gnd(gnd), .vdd(vdd), .B(_1513_), );
  NAND2X1 NAND2X1_344 (.Y(_2584_), .A(regs_18__3_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf84_), );
  NAND2X1 NAND2X1_345 (.Y(_2585_), .A(_2415__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_2584_), );
  OAI21X1 OAI21X1_1108 (.Y(_2586_), .A(_2585_), .gnd(gnd), .vdd(vdd), .B(_2583_), .C(raddr1_2_bF_buf5_), );
  OAI21X1 OAI21X1_1109 (.Y(_2587_), .A(_1414_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf83_), .C(raddr1_1_bF_buf0_), );
  AOI21X1 AOI21X1_142 (.Y(_2588_), .A(regs_20__3_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf82_), .C(_2587_), );
  AND2X2 AND2X2_5 (.Y(_2589_), .A(regs_22__3_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf81_), );
  OAI21X1 OAI21X1_1110 (.Y(_2590_), .A(_1316_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf80_), .C(_2415__bF_buf0), );
  OAI21X1 OAI21X1_1111 (.Y(_2591_), .A(_2590_), .gnd(gnd), .vdd(vdd), .B(_2589_), .C(_2399__bF_buf7), );
  OAI22X1 OAI22X1_6 (.Y(_2592_), .A(_2582_), .gnd(gnd), .vdd(vdd), .B(_2586_), .C(_2591_), .D(_2588_), );
  INVX1 INVX1_20 (.Y(_2593_), .A(regs_29__3_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_346 (.Y(_2594_), .A(regs_28__3_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf79_), );
  OAI21X1 OAI21X1_1112 (.Y(_2595_), .A(_2593_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf78_), .C(_2594_), );
  MUX2X1 MUX2X1_34 (.Y(_2596_), .A(_2595_), .gnd(gnd), .vdd(vdd), .B(regs_30__3_), .S(raddr1_1_bF_buf14_bF_buf1_), );
  NAND2X1 NAND2X1_347 (.Y(_2597_), .A(regs_26__3_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf77_), );
  OAI21X1 OAI21X1_1113 (.Y(_2598_), .A(_1149_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf76_), .C(_2597_), );
  INVX1 INVX1_21 (.Y(_2599_), .A(regs_25__3_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_348 (.Y(_2600_), .A(regs_24__3_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf75_), );
  OAI21X1 OAI21X1_1114 (.Y(_2601_), .A(_2599_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf74_), .C(_2600_), );
  MUX2X1 MUX2X1_35 (.Y(_2602_), .A(_2601_), .gnd(gnd), .vdd(vdd), .B(_2598_), .S(raddr1_1_bF_buf13_bF_buf1_), );
  MUX2X1 MUX2X1_36 (.Y(_2603_), .A(_2602_), .gnd(gnd), .vdd(vdd), .B(_2596_), .S(raddr1_2_bF_buf4_), );
  MUX2X1 MUX2X1_37 (.Y(_2604_), .A(_2603_), .gnd(gnd), .vdd(vdd), .B(_2592_), .S(_2398__bF_buf6), );
  MUX2X1 MUX2X1_38 (.Y(_5511__3_), .A(_2580_), .gnd(gnd), .vdd(vdd), .B(_2604_), .S(raddr1_4_bF_buf1_), );
  INVX1 INVX1_22 (.Y(_2605_), .A(regs_5__4_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1115 (.Y(_2606_), .A(_2605_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf73_), .C(raddr1_1_bF_buf12_bF_buf1_), );
  AOI21X1 AOI21X1_143 (.Y(_2607_), .A(regs_4__4_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf72_), .C(_2606_), );
  AND2X2 AND2X2_6 (.Y(_2608_), .A(regs_6__4_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf71_), );
  OAI21X1 OAI21X1_1116 (.Y(_2609_), .A(_2109_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf70_), .C(_2415__bF_buf8), );
  OAI21X1 OAI21X1_1117 (.Y(_2610_), .A(_2609_), .gnd(gnd), .vdd(vdd), .B(_2608_), .C(_2399__bF_buf6), );
  INVX1 INVX1_23 (.Y(_2611_), .A(regs_1__4_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1118 (.Y(_2612_), .A(_2611_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf69_), .C(raddr1_1_bF_buf11_bF_buf1_), );
  AOI21X1 AOI21X1_144 (.Y(_2613_), .A(regs_0__4_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf68_), .C(_2612_), );
  INVX1 INVX1_24 (.Y(_2614_), .A(regs_3__4_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_149 (.Y(_2615_), .A(raddr1_0_bF_buf67_), .gnd(gnd), .vdd(vdd), .B(_2614_), );
  NAND2X1 NAND2X1_349 (.Y(_2616_), .A(regs_2__4_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf66_), );
  NAND2X1 NAND2X1_350 (.Y(_2617_), .A(_2415__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_2616_), );
  OAI21X1 OAI21X1_1119 (.Y(_2618_), .A(_2617_), .gnd(gnd), .vdd(vdd), .B(_2615_), .C(raddr1_2_bF_buf3_), );
  OAI22X1 OAI22X1_7 (.Y(_2619_), .A(_2613_), .gnd(gnd), .vdd(vdd), .B(_2618_), .C(_2610_), .D(_2607_), );
  NAND2X1 NAND2X1_351 (.Y(_2620_), .A(regs_10__4_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf65_), );
  OAI21X1 OAI21X1_1120 (.Y(_2621_), .A(_1910_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf64_), .C(_2620_), );
  NAND2X1 NAND2X1_352 (.Y(_2622_), .A(regs_8__4_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf63_), );
  OAI21X1 OAI21X1_1121 (.Y(_2623_), .A(_2008_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf62_), .C(_2622_), );
  MUX2X1 MUX2X1_39 (.Y(_2624_), .A(_2623_), .gnd(gnd), .vdd(vdd), .B(_2621_), .S(raddr1_1_bF_buf10_bF_buf1_), );
  NAND2X1 NAND2X1_353 (.Y(_2625_), .A(regs_14__4_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf61_), );
  OAI21X1 OAI21X1_1122 (.Y(_2626_), .A(_1713_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf60_), .C(_2625_), );
  NAND2X1 NAND2X1_354 (.Y(_2627_), .A(regs_12__4_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf59_), );
  OAI21X1 OAI21X1_1123 (.Y(_2628_), .A(_1811_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf58_), .C(_2627_), );
  MUX2X1 MUX2X1_40 (.Y(_2629_), .A(_2628_), .gnd(gnd), .vdd(vdd), .B(_2626_), .S(raddr1_1_bF_buf9_bF_buf1_), );
  MUX2X1 MUX2X1_41 (.Y(_2630_), .A(_2629_), .gnd(gnd), .vdd(vdd), .B(_2624_), .S(_2399__bF_buf5), );
  MUX2X1 MUX2X1_42 (.Y(_2631_), .A(_2630_), .gnd(gnd), .vdd(vdd), .B(_2619_), .S(_2398__bF_buf5), );
  OAI21X1 OAI21X1_1124 (.Y(_2632_), .A(_1613_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf57_), .C(raddr1_1_bF_buf8_), );
  AOI21X1 AOI21X1_145 (.Y(_2633_), .A(regs_16__4_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf56_), .C(_2632_), );
  NOR2X1 NOR2X1_150 (.Y(_2634_), .A(raddr1_0_bF_buf55_), .gnd(gnd), .vdd(vdd), .B(_1515_), );
  NAND2X1 NAND2X1_355 (.Y(_2635_), .A(regs_18__4_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf54_), );
  NAND2X1 NAND2X1_356 (.Y(_2636_), .A(_2415__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_2635_), );
  OAI21X1 OAI21X1_1125 (.Y(_2637_), .A(_2636_), .gnd(gnd), .vdd(vdd), .B(_2634_), .C(raddr1_2_bF_buf2_), );
  OAI21X1 OAI21X1_1126 (.Y(_2638_), .A(_1416_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf53_), .C(raddr1_1_bF_buf7_), );
  AOI21X1 AOI21X1_146 (.Y(_2639_), .A(regs_20__4_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf52_), .C(_2638_), );
  AND2X2 AND2X2_7 (.Y(_2640_), .A(regs_22__4_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf51_), );
  OAI21X1 OAI21X1_1127 (.Y(_2641_), .A(_1318_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf50_), .C(_2415__bF_buf5), );
  OAI21X1 OAI21X1_1128 (.Y(_2642_), .A(_2641_), .gnd(gnd), .vdd(vdd), .B(_2640_), .C(_2399__bF_buf4), );
  OAI22X1 OAI22X1_8 (.Y(_2643_), .A(_2633_), .gnd(gnd), .vdd(vdd), .B(_2637_), .C(_2642_), .D(_2639_), );
  INVX1 INVX1_25 (.Y(_2644_), .A(regs_29__4_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_357 (.Y(_2645_), .A(regs_28__4_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf49_), );
  OAI21X1 OAI21X1_1129 (.Y(_2646_), .A(_2644_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf48_), .C(_2645_), );
  MUX2X1 MUX2X1_43 (.Y(_2647_), .A(_2646_), .gnd(gnd), .vdd(vdd), .B(regs_30__4_), .S(raddr1_1_bF_buf6_), );
  NAND2X1 NAND2X1_358 (.Y(_2648_), .A(regs_26__4_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf47_), );
  OAI21X1 OAI21X1_1130 (.Y(_2649_), .A(_1151_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf46_), .C(_2648_), );
  INVX1 INVX1_26 (.Y(_2650_), .A(regs_25__4_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_359 (.Y(_2651_), .A(regs_24__4_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf45_), );
  OAI21X1 OAI21X1_1131 (.Y(_2652_), .A(_2650_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf44_), .C(_2651_), );
  MUX2X1 MUX2X1_44 (.Y(_2653_), .A(_2652_), .gnd(gnd), .vdd(vdd), .B(_2649_), .S(raddr1_1_bF_buf5_), );
  MUX2X1 MUX2X1_45 (.Y(_2654_), .A(_2653_), .gnd(gnd), .vdd(vdd), .B(_2647_), .S(raddr1_2_bF_buf1_), );
  MUX2X1 MUX2X1_46 (.Y(_2655_), .A(_2654_), .gnd(gnd), .vdd(vdd), .B(_2643_), .S(_2398__bF_buf4), );
  MUX2X1 MUX2X1_47 (.Y(_5511__4_), .A(_2631_), .gnd(gnd), .vdd(vdd), .B(_2655_), .S(raddr1_4_bF_buf0_), );
  OAI21X1 OAI21X1_1132 (.Y(_2656_), .A(_1418_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf43_), .C(raddr1_1_bF_buf4_), );
  AOI21X1 AOI21X1_147 (.Y(_2657_), .A(regs_20__5_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf42_), .C(_2656_), );
  AND2X2 AND2X2_8 (.Y(_2658_), .A(regs_22__5_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf41_), );
  OAI21X1 OAI21X1_1133 (.Y(_2659_), .A(_1320_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf40_), .C(_2415__bF_buf4), );
  OAI21X1 OAI21X1_1134 (.Y(_2660_), .A(_2659_), .gnd(gnd), .vdd(vdd), .B(_2658_), .C(_2399__bF_buf3), );
  OAI21X1 OAI21X1_1135 (.Y(_2661_), .A(_1615_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf39_), .C(raddr1_1_bF_buf3_), );
  AOI21X1 AOI21X1_148 (.Y(_2662_), .A(regs_16__5_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf38_), .C(_2661_), );
  NOR2X1 NOR2X1_151 (.Y(_2663_), .A(raddr1_0_bF_buf37_), .gnd(gnd), .vdd(vdd), .B(_1517_), );
  NAND2X1 NAND2X1_360 (.Y(_2664_), .A(regs_18__5_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf36_), );
  NAND2X1 NAND2X1_361 (.Y(_2665_), .A(_2415__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_2664_), );
  OAI21X1 OAI21X1_1136 (.Y(_2666_), .A(_2665_), .gnd(gnd), .vdd(vdd), .B(_2663_), .C(raddr1_2_bF_buf0_), );
  OAI22X1 OAI22X1_9 (.Y(_2667_), .A(_2662_), .gnd(gnd), .vdd(vdd), .B(_2666_), .C(_2660_), .D(_2657_), );
  INVX1 INVX1_27 (.Y(_2668_), .A(regs_29__5_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_362 (.Y(_2669_), .A(regs_28__5_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf35_), );
  OAI21X1 OAI21X1_1137 (.Y(_2670_), .A(_2668_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf34_), .C(_2669_), );
  MUX2X1 MUX2X1_48 (.Y(_2671_), .A(_2670_), .gnd(gnd), .vdd(vdd), .B(regs_30__5_), .S(raddr1_1_bF_buf2_), );
  NAND2X1 NAND2X1_363 (.Y(_2672_), .A(regs_26__5_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf33_), );
  OAI21X1 OAI21X1_1138 (.Y(_2673_), .A(_1153_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf32_), .C(_2672_), );
  INVX1 INVX1_28 (.Y(_2674_), .A(regs_25__5_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_364 (.Y(_2675_), .A(regs_24__5_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf31_), );
  OAI21X1 OAI21X1_1139 (.Y(_2676_), .A(_2674_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf30_), .C(_2675_), );
  MUX2X1 MUX2X1_49 (.Y(_2677_), .A(_2676_), .gnd(gnd), .vdd(vdd), .B(_2673_), .S(raddr1_1_bF_buf1_), );
  MUX2X1 MUX2X1_50 (.Y(_2678_), .A(_2677_), .gnd(gnd), .vdd(vdd), .B(_2671_), .S(raddr1_2_bF_buf10_), );
  MUX2X1 MUX2X1_51 (.Y(_2679_), .A(_2678_), .gnd(gnd), .vdd(vdd), .B(_2667_), .S(_2398__bF_buf3), );
  NAND2X1 NAND2X1_365 (.Y(_2680_), .A(regs_6__5_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf29_), );
  OAI21X1 OAI21X1_1140 (.Y(_2681_), .A(_2111_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf28_), .C(_2680_), );
  INVX1 INVX1_29 (.Y(_2682_), .A(regs_5__5_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_366 (.Y(_2683_), .A(regs_4__5_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf27_), );
  OAI21X1 OAI21X1_1141 (.Y(_2684_), .A(_2682_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf26_), .C(_2683_), );
  MUX2X1 MUX2X1_52 (.Y(_2685_), .A(_2684_), .gnd(gnd), .vdd(vdd), .B(_2681_), .S(raddr1_1_bF_buf0_), );
  INVX1 INVX1_30 (.Y(_2686_), .A(regs_3__5_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_367 (.Y(_2687_), .A(regs_2__5_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf25_), );
  OAI21X1 OAI21X1_1142 (.Y(_2688_), .A(_2686_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf24_), .C(_2687_), );
  INVX1 INVX1_31 (.Y(_2689_), .A(regs_1__5_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_368 (.Y(_2690_), .A(regs_0__5_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf23_), );
  OAI21X1 OAI21X1_1143 (.Y(_2691_), .A(_2689_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf22_), .C(_2690_), );
  MUX2X1 MUX2X1_53 (.Y(_2692_), .A(_2691_), .gnd(gnd), .vdd(vdd), .B(_2688_), .S(raddr1_1_bF_buf14_bF_buf0_), );
  MUX2X1 MUX2X1_54 (.Y(_2693_), .A(_2692_), .gnd(gnd), .vdd(vdd), .B(_2685_), .S(raddr1_2_bF_buf9_), );
  NAND2X1 NAND2X1_369 (.Y(_2694_), .A(regs_14__5_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf21_), );
  OAI21X1 OAI21X1_1144 (.Y(_2695_), .A(_1715_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf20_), .C(_2694_), );
  NAND2X1 NAND2X1_370 (.Y(_2696_), .A(regs_12__5_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf19_), );
  OAI21X1 OAI21X1_1145 (.Y(_2697_), .A(_1813_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf18_), .C(_2696_), );
  MUX2X1 MUX2X1_55 (.Y(_2698_), .A(_2697_), .gnd(gnd), .vdd(vdd), .B(_2695_), .S(raddr1_1_bF_buf13_bF_buf0_), );
  NAND2X1 NAND2X1_371 (.Y(_2699_), .A(regs_10__5_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf17_), );
  OAI21X1 OAI21X1_1146 (.Y(_2700_), .A(_1912_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf16_), .C(_2699_), );
  NAND2X1 NAND2X1_372 (.Y(_2701_), .A(regs_8__5_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf15_), );
  OAI21X1 OAI21X1_1147 (.Y(_2702_), .A(_2010_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf14_), .C(_2701_), );
  MUX2X1 MUX2X1_56 (.Y(_2703_), .A(_2702_), .gnd(gnd), .vdd(vdd), .B(_2700_), .S(raddr1_1_bF_buf12_bF_buf0_), );
  MUX2X1 MUX2X1_57 (.Y(_2704_), .A(_2703_), .gnd(gnd), .vdd(vdd), .B(_2698_), .S(raddr1_2_bF_buf8_), );
  MUX2X1 MUX2X1_58 (.Y(_2705_), .A(_2704_), .gnd(gnd), .vdd(vdd), .B(_2693_), .S(_2398__bF_buf2), );
  MUX2X1 MUX2X1_59 (.Y(_5511__5_), .A(_2705_), .gnd(gnd), .vdd(vdd), .B(_2679_), .S(raddr1_4_bF_buf4_), );
  OAI21X1 OAI21X1_1148 (.Y(_2706_), .A(_1420_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf13_), .C(raddr1_1_bF_buf11_bF_buf0_), );
  AOI21X1 AOI21X1_149 (.Y(_2707_), .A(regs_20__6_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf12_), .C(_2706_), );
  AND2X2 AND2X2_9 (.Y(_2708_), .A(regs_22__6_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf11_), );
  OAI21X1 OAI21X1_1149 (.Y(_2709_), .A(_1322_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf10_), .C(_2415__bF_buf2), );
  OAI21X1 OAI21X1_1150 (.Y(_2710_), .A(_2709_), .gnd(gnd), .vdd(vdd), .B(_2708_), .C(_2399__bF_buf2), );
  OAI21X1 OAI21X1_1151 (.Y(_2711_), .A(_1617_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf9_), .C(raddr1_1_bF_buf10_bF_buf0_), );
  AOI21X1 AOI21X1_150 (.Y(_2712_), .A(regs_16__6_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf8_), .C(_2711_), );
  NOR2X1 NOR2X1_152 (.Y(_2713_), .A(raddr1_0_bF_buf7_), .gnd(gnd), .vdd(vdd), .B(_1519_), );
  NAND2X1 NAND2X1_373 (.Y(_2714_), .A(regs_18__6_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf6_), );
  NAND2X1 NAND2X1_374 (.Y(_2715_), .A(_2415__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_2714_), );
  OAI21X1 OAI21X1_1152 (.Y(_2716_), .A(_2715_), .gnd(gnd), .vdd(vdd), .B(_2713_), .C(raddr1_2_bF_buf7_), );
  OAI22X1 OAI22X1_10 (.Y(_2717_), .A(_2712_), .gnd(gnd), .vdd(vdd), .B(_2716_), .C(_2710_), .D(_2707_), );
  INVX1 INVX1_32 (.Y(_2718_), .A(regs_29__6_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_375 (.Y(_2719_), .A(regs_28__6_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf5_), );
  OAI21X1 OAI21X1_1153 (.Y(_2720_), .A(_2718_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf4_), .C(_2719_), );
  MUX2X1 MUX2X1_60 (.Y(_2721_), .A(_2720_), .gnd(gnd), .vdd(vdd), .B(regs_30__6_), .S(raddr1_1_bF_buf9_bF_buf0_), );
  NAND2X1 NAND2X1_376 (.Y(_2722_), .A(regs_26__6_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf3_), );
  OAI21X1 OAI21X1_1154 (.Y(_2723_), .A(_1155_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf2_), .C(_2722_), );
  INVX1 INVX1_33 (.Y(_2724_), .A(regs_25__6_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_377 (.Y(_2725_), .A(regs_24__6_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf1_), );
  OAI21X1 OAI21X1_1155 (.Y(_2726_), .A(_2724_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf0_), .C(_2725_), );
  MUX2X1 MUX2X1_61 (.Y(_2727_), .A(_2726_), .gnd(gnd), .vdd(vdd), .B(_2723_), .S(raddr1_1_bF_buf8_), );
  MUX2X1 MUX2X1_62 (.Y(_2728_), .A(_2727_), .gnd(gnd), .vdd(vdd), .B(_2721_), .S(raddr1_2_bF_buf6_), );
  MUX2X1 MUX2X1_63 (.Y(_2729_), .A(_2728_), .gnd(gnd), .vdd(vdd), .B(_2717_), .S(_2398__bF_buf1), );
  NAND2X1 NAND2X1_378 (.Y(_2730_), .A(regs_6__6_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf96_), );
  OAI21X1 OAI21X1_1156 (.Y(_2731_), .A(_2113_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf95_), .C(_2730_), );
  INVX1 INVX1_34 (.Y(_2732_), .A(regs_5__6_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_379 (.Y(_2733_), .A(regs_4__6_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf94_), );
  OAI21X1 OAI21X1_1157 (.Y(_2734_), .A(_2732_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf93_), .C(_2733_), );
  MUX2X1 MUX2X1_64 (.Y(_2735_), .A(_2734_), .gnd(gnd), .vdd(vdd), .B(_2731_), .S(raddr1_1_bF_buf7_), );
  INVX1 INVX1_35 (.Y(_2736_), .A(regs_3__6_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_380 (.Y(_2737_), .A(regs_2__6_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf92_), );
  OAI21X1 OAI21X1_1158 (.Y(_2738_), .A(_2736_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf91_), .C(_2737_), );
  INVX1 INVX1_36 (.Y(_2739_), .A(regs_1__6_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_381 (.Y(_2740_), .A(regs_0__6_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf90_), );
  OAI21X1 OAI21X1_1159 (.Y(_2741_), .A(_2739_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf89_), .C(_2740_), );
  MUX2X1 MUX2X1_65 (.Y(_2742_), .A(_2741_), .gnd(gnd), .vdd(vdd), .B(_2738_), .S(raddr1_1_bF_buf6_), );
  MUX2X1 MUX2X1_66 (.Y(_2743_), .A(_2742_), .gnd(gnd), .vdd(vdd), .B(_2735_), .S(raddr1_2_bF_buf5_), );
  NAND2X1 NAND2X1_382 (.Y(_2744_), .A(regs_14__6_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf88_), );
  OAI21X1 OAI21X1_1160 (.Y(_2745_), .A(_1717_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf87_), .C(_2744_), );
  NAND2X1 NAND2X1_383 (.Y(_2746_), .A(regs_12__6_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf86_), );
  OAI21X1 OAI21X1_1161 (.Y(_2747_), .A(_1815_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf85_), .C(_2746_), );
  MUX2X1 MUX2X1_67 (.Y(_2748_), .A(_2747_), .gnd(gnd), .vdd(vdd), .B(_2745_), .S(raddr1_1_bF_buf5_), );
  NAND2X1 NAND2X1_384 (.Y(_2749_), .A(regs_10__6_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf84_), );
  OAI21X1 OAI21X1_1162 (.Y(_2750_), .A(_1914_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf83_), .C(_2749_), );
  NAND2X1 NAND2X1_385 (.Y(_2751_), .A(regs_8__6_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf82_), );
  OAI21X1 OAI21X1_1163 (.Y(_2752_), .A(_2012_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf81_), .C(_2751_), );
  MUX2X1 MUX2X1_68 (.Y(_2753_), .A(_2752_), .gnd(gnd), .vdd(vdd), .B(_2750_), .S(raddr1_1_bF_buf4_), );
  MUX2X1 MUX2X1_69 (.Y(_2754_), .A(_2753_), .gnd(gnd), .vdd(vdd), .B(_2748_), .S(raddr1_2_bF_buf4_), );
  MUX2X1 MUX2X1_70 (.Y(_2755_), .A(_2754_), .gnd(gnd), .vdd(vdd), .B(_2743_), .S(_2398__bF_buf0), );
  MUX2X1 MUX2X1_71 (.Y(_5511__6_), .A(_2755_), .gnd(gnd), .vdd(vdd), .B(_2729_), .S(raddr1_4_bF_buf3_), );
  NAND2X1 NAND2X1_386 (.Y(_2756_), .A(regs_22__7_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf80_), );
  OAI21X1 OAI21X1_1164 (.Y(_2757_), .A(_1324_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf79_), .C(_2756_), );
  NAND2X1 NAND2X1_387 (.Y(_2758_), .A(regs_20__7_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf78_), );
  OAI21X1 OAI21X1_1165 (.Y(_2759_), .A(_1422_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf77_), .C(_2758_), );
  MUX2X1 MUX2X1_72 (.Y(_2760_), .A(_2759_), .gnd(gnd), .vdd(vdd), .B(_2757_), .S(raddr1_1_bF_buf3_), );
  NAND2X1 NAND2X1_388 (.Y(_2761_), .A(_2399__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_2760_), );
  NAND2X1 NAND2X1_389 (.Y(_2762_), .A(regs_18__7_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf76_), );
  OAI21X1 OAI21X1_1166 (.Y(_2763_), .A(_1521_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf75_), .C(_2762_), );
  NAND2X1 NAND2X1_390 (.Y(_2764_), .A(regs_16__7_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf74_), );
  OAI21X1 OAI21X1_1167 (.Y(_2765_), .A(_1619_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf73_), .C(_2764_), );
  MUX2X1 MUX2X1_73 (.Y(_2766_), .A(_2765_), .gnd(gnd), .vdd(vdd), .B(_2763_), .S(raddr1_1_bF_buf2_), );
  AOI21X1 AOI21X1_151 (.Y(_2767_), .A(raddr1_2_bF_buf3_), .gnd(gnd), .vdd(vdd), .B(_2766_), .C(_2398__bF_buf7), );
  OAI21X1 OAI21X1_1168 (.Y(_2768_), .A(_1157_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf72_), .C(raddr1_2_bF_buf2_), );
  AOI21X1 AOI21X1_152 (.Y(_2769_), .A(regs_26__7_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf71_), .C(_2768_), );
  OAI21X1 OAI21X1_1169 (.Y(_2770_), .A(regs_30__7_), .gnd(gnd), .vdd(vdd), .B(raddr1_2_bF_buf1_), .C(_2415__bF_buf0), );
  INVX1 INVX1_37 (.Y(_2771_), .A(regs_25__7_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1170 (.Y(_2772_), .A(_2771_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf70_), .C(raddr1_2_bF_buf0_), );
  AOI21X1 AOI21X1_153 (.Y(_2773_), .A(regs_24__7_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf69_), .C(_2772_), );
  INVX1 INVX1_38 (.Y(_2774_), .A(regs_29__7_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_153 (.Y(_2775_), .A(raddr1_0_bF_buf68_), .gnd(gnd), .vdd(vdd), .B(_2774_), );
  NAND2X1 NAND2X1_391 (.Y(_2776_), .A(regs_28__7_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf67_), );
  NAND2X1 NAND2X1_392 (.Y(_2777_), .A(_2399__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_2776_), );
  OAI21X1 OAI21X1_1171 (.Y(_2778_), .A(_2777_), .gnd(gnd), .vdd(vdd), .B(_2775_), .C(raddr1_1_bF_buf1_), );
  OAI22X1 OAI22X1_11 (.Y(_2779_), .A(_2769_), .gnd(gnd), .vdd(vdd), .B(_2770_), .C(_2778_), .D(_2773_), );
  AOI22X1 AOI22X1_3 (.Y(_2780_), .A(_2779_), .gnd(gnd), .vdd(vdd), .B(_2398__bF_buf6), .C(_2761_), .D(_2767_), );
  INVX1 INVX1_39 (.Y(_2781_), .A(regs_5__7_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1172 (.Y(_2782_), .A(_2781_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf66_), .C(raddr1_1_bF_buf0_), );
  AOI21X1 AOI21X1_154 (.Y(_2783_), .A(regs_4__7_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf65_), .C(_2782_), );
  AND2X2 AND2X2_10 (.Y(_2784_), .A(regs_6__7_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf64_), );
  OAI21X1 OAI21X1_1173 (.Y(_2785_), .A(_2115_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf63_), .C(_2415__bF_buf8), );
  OAI21X1 OAI21X1_1174 (.Y(_2786_), .A(_2785_), .gnd(gnd), .vdd(vdd), .B(_2784_), .C(_2399__bF_buf8), );
  INVX1 INVX1_40 (.Y(_2787_), .A(regs_1__7_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1175 (.Y(_2788_), .A(_2787_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf62_), .C(raddr1_1_bF_buf14_bF_buf3_), );
  AOI21X1 AOI21X1_155 (.Y(_2789_), .A(regs_0__7_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf61_), .C(_2788_), );
  INVX1 INVX1_41 (.Y(_2790_), .A(regs_3__7_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_154 (.Y(_2791_), .A(raddr1_0_bF_buf60_), .gnd(gnd), .vdd(vdd), .B(_2790_), );
  NAND2X1 NAND2X1_393 (.Y(_2792_), .A(regs_2__7_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf59_), );
  NAND2X1 NAND2X1_394 (.Y(_2793_), .A(_2415__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_2792_), );
  OAI21X1 OAI21X1_1176 (.Y(_2794_), .A(_2793_), .gnd(gnd), .vdd(vdd), .B(_2791_), .C(raddr1_2_bF_buf10_), );
  OAI22X1 OAI22X1_12 (.Y(_2795_), .A(_2789_), .gnd(gnd), .vdd(vdd), .B(_2794_), .C(_2786_), .D(_2783_), );
  NAND2X1 NAND2X1_395 (.Y(_2796_), .A(regs_10__7_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf58_), );
  OAI21X1 OAI21X1_1177 (.Y(_2797_), .A(_1916_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf57_), .C(_2796_), );
  NAND2X1 NAND2X1_396 (.Y(_2798_), .A(regs_8__7_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf56_), );
  OAI21X1 OAI21X1_1178 (.Y(_2799_), .A(_2014_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf55_), .C(_2798_), );
  MUX2X1 MUX2X1_74 (.Y(_2800_), .A(_2799_), .gnd(gnd), .vdd(vdd), .B(_2797_), .S(raddr1_1_bF_buf13_bF_buf3_), );
  NAND2X1 NAND2X1_397 (.Y(_2801_), .A(regs_14__7_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf54_), );
  OAI21X1 OAI21X1_1179 (.Y(_2802_), .A(_1719_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf53_), .C(_2801_), );
  NAND2X1 NAND2X1_398 (.Y(_2803_), .A(regs_12__7_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf52_), );
  OAI21X1 OAI21X1_1180 (.Y(_2804_), .A(_1817_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf51_), .C(_2803_), );
  MUX2X1 MUX2X1_75 (.Y(_2805_), .A(_2804_), .gnd(gnd), .vdd(vdd), .B(_2802_), .S(raddr1_1_bF_buf12_bF_buf3_), );
  MUX2X1 MUX2X1_76 (.Y(_2806_), .A(_2805_), .gnd(gnd), .vdd(vdd), .B(_2800_), .S(_2399__bF_buf7), );
  MUX2X1 MUX2X1_77 (.Y(_2807_), .A(_2806_), .gnd(gnd), .vdd(vdd), .B(_2795_), .S(_2398__bF_buf5), );
  MUX2X1 MUX2X1_78 (.Y(_5511__7_), .A(_2807_), .gnd(gnd), .vdd(vdd), .B(_2780_), .S(raddr1_4_bF_buf2_), );
  INVX1 INVX1_42 (.Y(_2808_), .A(regs_5__8_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1181 (.Y(_2809_), .A(_2808_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf50_), .C(raddr1_1_bF_buf11_bF_buf3_), );
  AOI21X1 AOI21X1_156 (.Y(_2810_), .A(regs_4__8_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf49_), .C(_2809_), );
  AND2X2 AND2X2_11 (.Y(_2811_), .A(regs_6__8_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf48_), );
  OAI21X1 OAI21X1_1182 (.Y(_2812_), .A(_2117_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf47_), .C(_2415__bF_buf6), );
  OAI21X1 OAI21X1_1183 (.Y(_2813_), .A(_2812_), .gnd(gnd), .vdd(vdd), .B(_2811_), .C(_2399__bF_buf6), );
  INVX1 INVX1_43 (.Y(_2814_), .A(regs_1__8_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1184 (.Y(_2815_), .A(_2814_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf46_), .C(raddr1_1_bF_buf10_bF_buf3_), );
  AOI21X1 AOI21X1_157 (.Y(_2816_), .A(regs_0__8_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf45_), .C(_2815_), );
  INVX1 INVX1_44 (.Y(_2817_), .A(regs_3__8_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_155 (.Y(_2818_), .A(raddr1_0_bF_buf44_), .gnd(gnd), .vdd(vdd), .B(_2817_), );
  NAND2X1 NAND2X1_399 (.Y(_2819_), .A(regs_2__8_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf43_), );
  NAND2X1 NAND2X1_400 (.Y(_2820_), .A(_2415__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_2819_), );
  OAI21X1 OAI21X1_1185 (.Y(_2821_), .A(_2820_), .gnd(gnd), .vdd(vdd), .B(_2818_), .C(raddr1_2_bF_buf9_), );
  OAI22X1 OAI22X1_13 (.Y(_2822_), .A(_2816_), .gnd(gnd), .vdd(vdd), .B(_2821_), .C(_2813_), .D(_2810_), );
  NAND2X1 NAND2X1_401 (.Y(_2823_), .A(regs_10__8_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf42_), );
  OAI21X1 OAI21X1_1186 (.Y(_2824_), .A(_1918_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf41_), .C(_2823_), );
  NAND2X1 NAND2X1_402 (.Y(_2825_), .A(regs_8__8_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf40_), );
  OAI21X1 OAI21X1_1187 (.Y(_2826_), .A(_2016_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf39_), .C(_2825_), );
  MUX2X1 MUX2X1_79 (.Y(_2827_), .A(_2826_), .gnd(gnd), .vdd(vdd), .B(_2824_), .S(raddr1_1_bF_buf9_bF_buf3_), );
  NAND2X1 NAND2X1_403 (.Y(_2828_), .A(regs_14__8_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf38_), );
  OAI21X1 OAI21X1_1188 (.Y(_2829_), .A(_1721_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf37_), .C(_2828_), );
  NAND2X1 NAND2X1_404 (.Y(_2830_), .A(regs_12__8_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf36_), );
  OAI21X1 OAI21X1_1189 (.Y(_2831_), .A(_1819_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf35_), .C(_2830_), );
  MUX2X1 MUX2X1_80 (.Y(_2832_), .A(_2831_), .gnd(gnd), .vdd(vdd), .B(_2829_), .S(raddr1_1_bF_buf8_), );
  MUX2X1 MUX2X1_81 (.Y(_2833_), .A(_2832_), .gnd(gnd), .vdd(vdd), .B(_2827_), .S(_2399__bF_buf5), );
  MUX2X1 MUX2X1_82 (.Y(_2834_), .A(_2833_), .gnd(gnd), .vdd(vdd), .B(_2822_), .S(_2398__bF_buf4), );
  OAI21X1 OAI21X1_1190 (.Y(_2835_), .A(_1621_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf34_), .C(raddr1_1_bF_buf7_), );
  AOI21X1 AOI21X1_158 (.Y(_2836_), .A(regs_16__8_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf33_), .C(_2835_), );
  NOR2X1 NOR2X1_156 (.Y(_2837_), .A(raddr1_0_bF_buf32_), .gnd(gnd), .vdd(vdd), .B(_1523_), );
  NAND2X1 NAND2X1_405 (.Y(_2838_), .A(regs_18__8_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf31_), );
  NAND2X1 NAND2X1_406 (.Y(_2839_), .A(_2415__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_2838_), );
  OAI21X1 OAI21X1_1191 (.Y(_2840_), .A(_2839_), .gnd(gnd), .vdd(vdd), .B(_2837_), .C(raddr1_2_bF_buf8_), );
  OAI21X1 OAI21X1_1192 (.Y(_2841_), .A(_1424_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf30_), .C(raddr1_1_bF_buf6_), );
  AOI21X1 AOI21X1_159 (.Y(_2842_), .A(regs_20__8_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf29_), .C(_2841_), );
  AND2X2 AND2X2_12 (.Y(_2843_), .A(regs_22__8_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf28_), );
  OAI21X1 OAI21X1_1193 (.Y(_2844_), .A(_1326_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf27_), .C(_2415__bF_buf3), );
  OAI21X1 OAI21X1_1194 (.Y(_2845_), .A(_2844_), .gnd(gnd), .vdd(vdd), .B(_2843_), .C(_2399__bF_buf4), );
  OAI22X1 OAI22X1_14 (.Y(_2846_), .A(_2836_), .gnd(gnd), .vdd(vdd), .B(_2840_), .C(_2845_), .D(_2842_), );
  INVX1 INVX1_45 (.Y(_2847_), .A(regs_29__8_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_407 (.Y(_2848_), .A(regs_28__8_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf26_), );
  OAI21X1 OAI21X1_1195 (.Y(_2849_), .A(_2847_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf25_), .C(_2848_), );
  MUX2X1 MUX2X1_83 (.Y(_2850_), .A(_2849_), .gnd(gnd), .vdd(vdd), .B(regs_30__8_), .S(raddr1_1_bF_buf5_), );
  NAND2X1 NAND2X1_408 (.Y(_2851_), .A(regs_26__8_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf24_), );
  OAI21X1 OAI21X1_1196 (.Y(_2852_), .A(_1159_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf23_), .C(_2851_), );
  INVX1 INVX1_46 (.Y(_2853_), .A(regs_25__8_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_409 (.Y(_2854_), .A(regs_24__8_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf22_), );
  OAI21X1 OAI21X1_1197 (.Y(_2855_), .A(_2853_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf21_), .C(_2854_), );
  MUX2X1 MUX2X1_84 (.Y(_2856_), .A(_2855_), .gnd(gnd), .vdd(vdd), .B(_2852_), .S(raddr1_1_bF_buf4_), );
  MUX2X1 MUX2X1_85 (.Y(_2857_), .A(_2856_), .gnd(gnd), .vdd(vdd), .B(_2850_), .S(raddr1_2_bF_buf7_), );
  MUX2X1 MUX2X1_86 (.Y(_2858_), .A(_2857_), .gnd(gnd), .vdd(vdd), .B(_2846_), .S(_2398__bF_buf3), );
  MUX2X1 MUX2X1_87 (.Y(_5511__8_), .A(_2834_), .gnd(gnd), .vdd(vdd), .B(_2858_), .S(raddr1_4_bF_buf1_), );
  NAND2X1 NAND2X1_410 (.Y(_2859_), .A(regs_22__9_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf20_), );
  OAI21X1 OAI21X1_1198 (.Y(_2860_), .A(_1328_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf19_), .C(_2859_), );
  NAND2X1 NAND2X1_411 (.Y(_2861_), .A(regs_20__9_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf18_), );
  OAI21X1 OAI21X1_1199 (.Y(_2862_), .A(_1426_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf17_), .C(_2861_), );
  MUX2X1 MUX2X1_88 (.Y(_2863_), .A(_2862_), .gnd(gnd), .vdd(vdd), .B(_2860_), .S(raddr1_1_bF_buf3_), );
  NAND2X1 NAND2X1_412 (.Y(_2864_), .A(_2399__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_2863_), );
  NAND2X1 NAND2X1_413 (.Y(_2865_), .A(regs_18__9_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf16_), );
  OAI21X1 OAI21X1_1200 (.Y(_2866_), .A(_1525_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf15_), .C(_2865_), );
  NAND2X1 NAND2X1_414 (.Y(_2867_), .A(regs_16__9_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf14_), );
  OAI21X1 OAI21X1_1201 (.Y(_2868_), .A(_1623_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf13_), .C(_2867_), );
  MUX2X1 MUX2X1_89 (.Y(_2869_), .A(_2868_), .gnd(gnd), .vdd(vdd), .B(_2866_), .S(raddr1_1_bF_buf2_), );
  AOI21X1 AOI21X1_160 (.Y(_2870_), .A(raddr1_2_bF_buf6_), .gnd(gnd), .vdd(vdd), .B(_2869_), .C(_2398__bF_buf2), );
  OAI21X1 OAI21X1_1202 (.Y(_2871_), .A(_1161_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf12_), .C(raddr1_2_bF_buf5_), );
  AOI21X1 AOI21X1_161 (.Y(_2872_), .A(regs_26__9_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf11_), .C(_2871_), );
  OAI21X1 OAI21X1_1203 (.Y(_2873_), .A(regs_30__9_), .gnd(gnd), .vdd(vdd), .B(raddr1_2_bF_buf4_), .C(_2415__bF_buf2), );
  INVX1 INVX1_47 (.Y(_2874_), .A(regs_25__9_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1204 (.Y(_2875_), .A(_2874_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf10_), .C(raddr1_2_bF_buf3_), );
  AOI21X1 AOI21X1_162 (.Y(_2876_), .A(regs_24__9_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf9_), .C(_2875_), );
  INVX1 INVX1_48 (.Y(_2877_), .A(regs_29__9_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_157 (.Y(_2878_), .A(raddr1_0_bF_buf8_), .gnd(gnd), .vdd(vdd), .B(_2877_), );
  NAND2X1 NAND2X1_415 (.Y(_2879_), .A(regs_28__9_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf7_), );
  NAND2X1 NAND2X1_416 (.Y(_2880_), .A(_2399__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_2879_), );
  OAI21X1 OAI21X1_1205 (.Y(_2881_), .A(_2880_), .gnd(gnd), .vdd(vdd), .B(_2878_), .C(raddr1_1_bF_buf1_), );
  OAI22X1 OAI22X1_15 (.Y(_2882_), .A(_2872_), .gnd(gnd), .vdd(vdd), .B(_2873_), .C(_2881_), .D(_2876_), );
  AOI22X1 AOI22X1_4 (.Y(_2883_), .A(_2882_), .gnd(gnd), .vdd(vdd), .B(_2398__bF_buf1), .C(_2864_), .D(_2870_), );
  NAND2X1 NAND2X1_417 (.Y(_2884_), .A(regs_6__9_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf6_), );
  OAI21X1 OAI21X1_1206 (.Y(_2885_), .A(_2119_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf5_), .C(_2884_), );
  INVX1 INVX1_49 (.Y(_2886_), .A(regs_5__9_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_418 (.Y(_2887_), .A(regs_4__9_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf4_), );
  OAI21X1 OAI21X1_1207 (.Y(_2888_), .A(_2886_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf3_), .C(_2887_), );
  MUX2X1 MUX2X1_90 (.Y(_2889_), .A(_2888_), .gnd(gnd), .vdd(vdd), .B(_2885_), .S(raddr1_1_bF_buf0_), );
  INVX1 INVX1_50 (.Y(_2890_), .A(regs_3__9_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_419 (.Y(_2891_), .A(regs_2__9_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf2_), );
  OAI21X1 OAI21X1_1208 (.Y(_2892_), .A(_2890_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf1_), .C(_2891_), );
  INVX1 INVX1_51 (.Y(_2893_), .A(regs_1__9_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_420 (.Y(_2894_), .A(regs_0__9_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf0_), );
  OAI21X1 OAI21X1_1209 (.Y(_2895_), .A(_2893_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf96_), .C(_2894_), );
  MUX2X1 MUX2X1_91 (.Y(_2896_), .A(_2895_), .gnd(gnd), .vdd(vdd), .B(_2892_), .S(raddr1_1_bF_buf14_bF_buf2_), );
  MUX2X1 MUX2X1_92 (.Y(_2897_), .A(_2896_), .gnd(gnd), .vdd(vdd), .B(_2889_), .S(raddr1_2_bF_buf2_), );
  NAND2X1 NAND2X1_421 (.Y(_2898_), .A(regs_14__9_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf95_), );
  OAI21X1 OAI21X1_1210 (.Y(_2899_), .A(_1723_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf94_), .C(_2898_), );
  NAND2X1 NAND2X1_422 (.Y(_2900_), .A(regs_12__9_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf93_), );
  OAI21X1 OAI21X1_1211 (.Y(_2901_), .A(_1821_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf92_), .C(_2900_), );
  MUX2X1 MUX2X1_93 (.Y(_2902_), .A(_2901_), .gnd(gnd), .vdd(vdd), .B(_2899_), .S(raddr1_1_bF_buf13_bF_buf2_), );
  NAND2X1 NAND2X1_423 (.Y(_2903_), .A(regs_10__9_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf91_), );
  OAI21X1 OAI21X1_1212 (.Y(_2904_), .A(_1920_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf90_), .C(_2903_), );
  NAND2X1 NAND2X1_424 (.Y(_2905_), .A(regs_8__9_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf89_), );
  OAI21X1 OAI21X1_1213 (.Y(_2906_), .A(_2018_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf88_), .C(_2905_), );
  MUX2X1 MUX2X1_94 (.Y(_2907_), .A(_2906_), .gnd(gnd), .vdd(vdd), .B(_2904_), .S(raddr1_1_bF_buf12_bF_buf2_), );
  MUX2X1 MUX2X1_95 (.Y(_2908_), .A(_2907_), .gnd(gnd), .vdd(vdd), .B(_2902_), .S(raddr1_2_bF_buf1_), );
  MUX2X1 MUX2X1_96 (.Y(_2909_), .A(_2908_), .gnd(gnd), .vdd(vdd), .B(_2897_), .S(_2398__bF_buf0), );
  MUX2X1 MUX2X1_97 (.Y(_5511__9_), .A(_2909_), .gnd(gnd), .vdd(vdd), .B(_2883_), .S(raddr1_4_bF_buf0_), );
  NAND2X1 NAND2X1_425 (.Y(_2910_), .A(regs_22__10_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf87_), );
  OAI21X1 OAI21X1_1214 (.Y(_2911_), .A(_1330_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf86_), .C(_2910_), );
  NAND2X1 NAND2X1_426 (.Y(_2912_), .A(regs_20__10_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf85_), );
  OAI21X1 OAI21X1_1215 (.Y(_2913_), .A(_1428_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf84_), .C(_2912_), );
  MUX2X1 MUX2X1_98 (.Y(_2914_), .A(_2913_), .gnd(gnd), .vdd(vdd), .B(_2911_), .S(raddr1_1_bF_buf11_bF_buf2_), );
  NAND2X1 NAND2X1_427 (.Y(_2915_), .A(_2399__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_2914_), );
  NAND2X1 NAND2X1_428 (.Y(_2916_), .A(regs_18__10_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf83_), );
  OAI21X1 OAI21X1_1216 (.Y(_2917_), .A(_1527_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf82_), .C(_2916_), );
  NAND2X1 NAND2X1_429 (.Y(_2918_), .A(regs_16__10_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf81_), );
  OAI21X1 OAI21X1_1217 (.Y(_2919_), .A(_1625_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf80_), .C(_2918_), );
  MUX2X1 MUX2X1_99 (.Y(_2920_), .A(_2919_), .gnd(gnd), .vdd(vdd), .B(_2917_), .S(raddr1_1_bF_buf10_bF_buf2_), );
  AOI21X1 AOI21X1_163 (.Y(_2921_), .A(raddr1_2_bF_buf0_), .gnd(gnd), .vdd(vdd), .B(_2920_), .C(_2398__bF_buf7), );
  OAI21X1 OAI21X1_1218 (.Y(_2922_), .A(_1163_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf79_), .C(raddr1_2_bF_buf10_), );
  AOI21X1 AOI21X1_164 (.Y(_2923_), .A(regs_26__10_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf78_), .C(_2922_), );
  OAI21X1 OAI21X1_1219 (.Y(_2924_), .A(regs_30__10_), .gnd(gnd), .vdd(vdd), .B(raddr1_2_bF_buf9_), .C(_2415__bF_buf1), );
  INVX1 INVX1_52 (.Y(_2925_), .A(regs_25__10_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1220 (.Y(_2926_), .A(_2925_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf77_), .C(raddr1_2_bF_buf8_), );
  AOI21X1 AOI21X1_165 (.Y(_2927_), .A(regs_24__10_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf76_), .C(_2926_), );
  INVX1 INVX1_53 (.Y(_2928_), .A(regs_29__10_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_158 (.Y(_2929_), .A(raddr1_0_bF_buf75_), .gnd(gnd), .vdd(vdd), .B(_2928_), );
  NAND2X1 NAND2X1_430 (.Y(_2930_), .A(regs_28__10_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf74_), );
  NAND2X1 NAND2X1_431 (.Y(_2931_), .A(_2399__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_2930_), );
  OAI21X1 OAI21X1_1221 (.Y(_2932_), .A(_2931_), .gnd(gnd), .vdd(vdd), .B(_2929_), .C(raddr1_1_bF_buf9_bF_buf2_), );
  OAI22X1 OAI22X1_16 (.Y(_2933_), .A(_2923_), .gnd(gnd), .vdd(vdd), .B(_2924_), .C(_2932_), .D(_2927_), );
  AOI22X1 AOI22X1_5 (.Y(_2934_), .A(_2933_), .gnd(gnd), .vdd(vdd), .B(_2398__bF_buf6), .C(_2915_), .D(_2921_), );
  INVX1 INVX1_54 (.Y(_2935_), .A(regs_5__10_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1222 (.Y(_2936_), .A(_2935_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf73_), .C(raddr1_1_bF_buf8_), );
  AOI21X1 AOI21X1_166 (.Y(_2937_), .A(regs_4__10_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf72_), .C(_2936_), );
  AND2X2 AND2X2_13 (.Y(_2938_), .A(regs_6__10_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf71_), );
  OAI21X1 OAI21X1_1223 (.Y(_2939_), .A(_2121_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf70_), .C(_2415__bF_buf0), );
  OAI21X1 OAI21X1_1224 (.Y(_2940_), .A(_2939_), .gnd(gnd), .vdd(vdd), .B(_2938_), .C(_2399__bF_buf8), );
  INVX1 INVX1_55 (.Y(_2941_), .A(regs_1__10_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1225 (.Y(_2942_), .A(_2941_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf69_), .C(raddr1_1_bF_buf7_), );
  AOI21X1 AOI21X1_167 (.Y(_2943_), .A(regs_0__10_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf68_), .C(_2942_), );
  INVX1 INVX1_56 (.Y(_2944_), .A(regs_3__10_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_159 (.Y(_2945_), .A(raddr1_0_bF_buf67_), .gnd(gnd), .vdd(vdd), .B(_2944_), );
  NAND2X1 NAND2X1_432 (.Y(_2946_), .A(regs_2__10_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf66_), );
  NAND2X1 NAND2X1_433 (.Y(_2947_), .A(_2415__bF_buf8), .gnd(gnd), .vdd(vdd), .B(_2946_), );
  OAI21X1 OAI21X1_1226 (.Y(_2948_), .A(_2947_), .gnd(gnd), .vdd(vdd), .B(_2945_), .C(raddr1_2_bF_buf7_), );
  OAI22X1 OAI22X1_17 (.Y(_2949_), .A(_2943_), .gnd(gnd), .vdd(vdd), .B(_2948_), .C(_2940_), .D(_2937_), );
  NAND2X1 NAND2X1_434 (.Y(_2950_), .A(regs_10__10_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf65_), );
  OAI21X1 OAI21X1_1227 (.Y(_2951_), .A(_1922_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf64_), .C(_2950_), );
  NAND2X1 NAND2X1_435 (.Y(_2952_), .A(regs_8__10_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf63_), );
  OAI21X1 OAI21X1_1228 (.Y(_2953_), .A(_2020_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf62_), .C(_2952_), );
  MUX2X1 MUX2X1_100 (.Y(_2954_), .A(_2953_), .gnd(gnd), .vdd(vdd), .B(_2951_), .S(raddr1_1_bF_buf6_), );
  NAND2X1 NAND2X1_436 (.Y(_2955_), .A(regs_14__10_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf61_), );
  OAI21X1 OAI21X1_1229 (.Y(_2956_), .A(_1725_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf60_), .C(_2955_), );
  NAND2X1 NAND2X1_437 (.Y(_2957_), .A(regs_12__10_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf59_), );
  OAI21X1 OAI21X1_1230 (.Y(_2958_), .A(_1823_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf58_), .C(_2957_), );
  MUX2X1 MUX2X1_101 (.Y(_2959_), .A(_2958_), .gnd(gnd), .vdd(vdd), .B(_2956_), .S(raddr1_1_bF_buf5_), );
  MUX2X1 MUX2X1_102 (.Y(_2960_), .A(_2959_), .gnd(gnd), .vdd(vdd), .B(_2954_), .S(_2399__bF_buf7), );
  MUX2X1 MUX2X1_103 (.Y(_2961_), .A(_2960_), .gnd(gnd), .vdd(vdd), .B(_2949_), .S(_2398__bF_buf5), );
  MUX2X1 MUX2X1_104 (.Y(_5511__10_), .A(_2961_), .gnd(gnd), .vdd(vdd), .B(_2934_), .S(raddr1_4_bF_buf4_), );
  INVX1 INVX1_57 (.Y(_2962_), .A(regs_5__11_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1231 (.Y(_2963_), .A(_2962_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf57_), .C(raddr1_1_bF_buf4_), );
  AOI21X1 AOI21X1_168 (.Y(_2964_), .A(regs_4__11_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf56_), .C(_2963_), );
  AND2X2 AND2X2_14 (.Y(_2965_), .A(regs_6__11_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf55_), );
  OAI21X1 OAI21X1_1232 (.Y(_2966_), .A(_2123_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf54_), .C(_2415__bF_buf7), );
  OAI21X1 OAI21X1_1233 (.Y(_2967_), .A(_2966_), .gnd(gnd), .vdd(vdd), .B(_2965_), .C(_2399__bF_buf6), );
  INVX1 INVX1_58 (.Y(_2968_), .A(regs_1__11_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1234 (.Y(_2969_), .A(_2968_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf53_), .C(raddr1_1_bF_buf3_), );
  AOI21X1 AOI21X1_169 (.Y(_2970_), .A(regs_0__11_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf52_), .C(_2969_), );
  INVX1 INVX1_59 (.Y(_2971_), .A(regs_3__11_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_160 (.Y(_2972_), .A(raddr1_0_bF_buf51_), .gnd(gnd), .vdd(vdd), .B(_2971_), );
  NAND2X1 NAND2X1_438 (.Y(_2973_), .A(regs_2__11_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf50_), );
  NAND2X1 NAND2X1_439 (.Y(_2974_), .A(_2415__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_2973_), );
  OAI21X1 OAI21X1_1235 (.Y(_2975_), .A(_2974_), .gnd(gnd), .vdd(vdd), .B(_2972_), .C(raddr1_2_bF_buf6_), );
  OAI22X1 OAI22X1_18 (.Y(_2976_), .A(_2970_), .gnd(gnd), .vdd(vdd), .B(_2975_), .C(_2967_), .D(_2964_), );
  NAND2X1 NAND2X1_440 (.Y(_2977_), .A(regs_10__11_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf49_), );
  OAI21X1 OAI21X1_1236 (.Y(_2978_), .A(_1924_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf48_), .C(_2977_), );
  NAND2X1 NAND2X1_441 (.Y(_2979_), .A(regs_8__11_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf47_), );
  OAI21X1 OAI21X1_1237 (.Y(_2980_), .A(_2022_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf46_), .C(_2979_), );
  MUX2X1 MUX2X1_105 (.Y(_2981_), .A(_2980_), .gnd(gnd), .vdd(vdd), .B(_2978_), .S(raddr1_1_bF_buf2_), );
  NAND2X1 NAND2X1_442 (.Y(_2982_), .A(regs_14__11_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf45_), );
  OAI21X1 OAI21X1_1238 (.Y(_2983_), .A(_1727_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf44_), .C(_2982_), );
  NAND2X1 NAND2X1_443 (.Y(_2984_), .A(regs_12__11_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf43_), );
  OAI21X1 OAI21X1_1239 (.Y(_2985_), .A(_1825_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf42_), .C(_2984_), );
  MUX2X1 MUX2X1_106 (.Y(_2986_), .A(_2985_), .gnd(gnd), .vdd(vdd), .B(_2983_), .S(raddr1_1_bF_buf1_), );
  MUX2X1 MUX2X1_107 (.Y(_2987_), .A(_2986_), .gnd(gnd), .vdd(vdd), .B(_2981_), .S(_2399__bF_buf5), );
  MUX2X1 MUX2X1_108 (.Y(_2988_), .A(_2987_), .gnd(gnd), .vdd(vdd), .B(_2976_), .S(_2398__bF_buf4), );
  OAI21X1 OAI21X1_1240 (.Y(_2989_), .A(_1627_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf41_), .C(raddr1_1_bF_buf0_), );
  AOI21X1 AOI21X1_170 (.Y(_2990_), .A(regs_16__11_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf40_), .C(_2989_), );
  NOR2X1 NOR2X1_161 (.Y(_2991_), .A(raddr1_0_bF_buf39_), .gnd(gnd), .vdd(vdd), .B(_1529_), );
  NAND2X1 NAND2X1_444 (.Y(_2992_), .A(regs_18__11_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf38_), );
  NAND2X1 NAND2X1_445 (.Y(_2993_), .A(_2415__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_2992_), );
  OAI21X1 OAI21X1_1241 (.Y(_2994_), .A(_2993_), .gnd(gnd), .vdd(vdd), .B(_2991_), .C(raddr1_2_bF_buf5_), );
  OAI21X1 OAI21X1_1242 (.Y(_2995_), .A(_1430_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf37_), .C(raddr1_1_bF_buf14_bF_buf1_), );
  AOI21X1 AOI21X1_171 (.Y(_2996_), .A(regs_20__11_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf36_), .C(_2995_), );
  AND2X2 AND2X2_15 (.Y(_2997_), .A(regs_22__11_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf35_), );
  OAI21X1 OAI21X1_1243 (.Y(_2998_), .A(_1332_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf34_), .C(_2415__bF_buf4), );
  OAI21X1 OAI21X1_1244 (.Y(_2999_), .A(_2998_), .gnd(gnd), .vdd(vdd), .B(_2997_), .C(_2399__bF_buf4), );
  OAI22X1 OAI22X1_19 (.Y(_3000_), .A(_2990_), .gnd(gnd), .vdd(vdd), .B(_2994_), .C(_2999_), .D(_2996_), );
  INVX1 INVX1_60 (.Y(_3001_), .A(regs_29__11_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_446 (.Y(_3002_), .A(regs_28__11_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf33_), );
  OAI21X1 OAI21X1_1245 (.Y(_3003_), .A(_3001_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf32_), .C(_3002_), );
  MUX2X1 MUX2X1_109 (.Y(_3004_), .A(_3003_), .gnd(gnd), .vdd(vdd), .B(regs_30__11_), .S(raddr1_1_bF_buf13_bF_buf1_), );
  NAND2X1 NAND2X1_447 (.Y(_3005_), .A(regs_26__11_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf31_), );
  OAI21X1 OAI21X1_1246 (.Y(_3006_), .A(_1165_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf30_), .C(_3005_), );
  INVX1 INVX1_61 (.Y(_3007_), .A(regs_25__11_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_448 (.Y(_3008_), .A(regs_24__11_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf29_), );
  OAI21X1 OAI21X1_1247 (.Y(_3009_), .A(_3007_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf28_), .C(_3008_), );
  MUX2X1 MUX2X1_110 (.Y(_3010_), .A(_3009_), .gnd(gnd), .vdd(vdd), .B(_3006_), .S(raddr1_1_bF_buf12_bF_buf1_), );
  MUX2X1 MUX2X1_111 (.Y(_3011_), .A(_3010_), .gnd(gnd), .vdd(vdd), .B(_3004_), .S(raddr1_2_bF_buf4_), );
  MUX2X1 MUX2X1_112 (.Y(_3012_), .A(_3011_), .gnd(gnd), .vdd(vdd), .B(_3000_), .S(_2398__bF_buf3), );
  MUX2X1 MUX2X1_113 (.Y(_5511__11_), .A(_2988_), .gnd(gnd), .vdd(vdd), .B(_3012_), .S(raddr1_4_bF_buf3_), );
  INVX1 INVX1_62 (.Y(_3013_), .A(regs_5__12_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1248 (.Y(_3014_), .A(_3013_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf27_), .C(raddr1_1_bF_buf11_bF_buf1_), );
  AOI21X1 AOI21X1_172 (.Y(_3015_), .A(regs_4__12_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf26_), .C(_3014_), );
  AND2X2 AND2X2_16 (.Y(_3016_), .A(regs_6__12_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf25_), );
  OAI21X1 OAI21X1_1249 (.Y(_3017_), .A(_2125_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf24_), .C(_2415__bF_buf3), );
  OAI21X1 OAI21X1_1250 (.Y(_3018_), .A(_3017_), .gnd(gnd), .vdd(vdd), .B(_3016_), .C(_2399__bF_buf3), );
  INVX1 INVX1_63 (.Y(_3019_), .A(regs_1__12_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1251 (.Y(_3020_), .A(_3019_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf23_), .C(raddr1_1_bF_buf10_bF_buf1_), );
  AOI21X1 AOI21X1_173 (.Y(_3021_), .A(regs_0__12_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf22_), .C(_3020_), );
  INVX1 INVX1_64 (.Y(_3022_), .A(regs_3__12_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_162 (.Y(_3023_), .A(raddr1_0_bF_buf21_), .gnd(gnd), .vdd(vdd), .B(_3022_), );
  NAND2X1 NAND2X1_449 (.Y(_3024_), .A(regs_2__12_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf20_), );
  NAND2X1 NAND2X1_450 (.Y(_3025_), .A(_2415__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_3024_), );
  OAI21X1 OAI21X1_1252 (.Y(_3026_), .A(_3025_), .gnd(gnd), .vdd(vdd), .B(_3023_), .C(raddr1_2_bF_buf3_), );
  OAI22X1 OAI22X1_20 (.Y(_3027_), .A(_3021_), .gnd(gnd), .vdd(vdd), .B(_3026_), .C(_3018_), .D(_3015_), );
  NAND2X1 NAND2X1_451 (.Y(_3028_), .A(regs_10__12_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf19_), );
  OAI21X1 OAI21X1_1253 (.Y(_3029_), .A(_1926_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf18_), .C(_3028_), );
  NAND2X1 NAND2X1_452 (.Y(_3030_), .A(regs_8__12_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf17_), );
  OAI21X1 OAI21X1_1254 (.Y(_3031_), .A(_2024_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf16_), .C(_3030_), );
  MUX2X1 MUX2X1_114 (.Y(_3032_), .A(_3031_), .gnd(gnd), .vdd(vdd), .B(_3029_), .S(raddr1_1_bF_buf9_bF_buf1_), );
  NAND2X1 NAND2X1_453 (.Y(_3033_), .A(regs_14__12_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf15_), );
  OAI21X1 OAI21X1_1255 (.Y(_3034_), .A(_1729_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf14_), .C(_3033_), );
  NAND2X1 NAND2X1_454 (.Y(_3035_), .A(regs_12__12_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf13_), );
  OAI21X1 OAI21X1_1256 (.Y(_3036_), .A(_1827_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf12_), .C(_3035_), );
  MUX2X1 MUX2X1_115 (.Y(_3037_), .A(_3036_), .gnd(gnd), .vdd(vdd), .B(_3034_), .S(raddr1_1_bF_buf8_), );
  MUX2X1 MUX2X1_116 (.Y(_3038_), .A(_3037_), .gnd(gnd), .vdd(vdd), .B(_3032_), .S(_2399__bF_buf2), );
  MUX2X1 MUX2X1_117 (.Y(_3039_), .A(_3038_), .gnd(gnd), .vdd(vdd), .B(_3027_), .S(_2398__bF_buf2), );
  OAI21X1 OAI21X1_1257 (.Y(_3040_), .A(_1629_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf11_), .C(raddr1_1_bF_buf7_), );
  AOI21X1 AOI21X1_174 (.Y(_3041_), .A(regs_16__12_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf10_), .C(_3040_), );
  NOR2X1 NOR2X1_163 (.Y(_3042_), .A(raddr1_0_bF_buf9_), .gnd(gnd), .vdd(vdd), .B(_1531_), );
  NAND2X1 NAND2X1_455 (.Y(_3043_), .A(regs_18__12_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf8_), );
  NAND2X1 NAND2X1_456 (.Y(_3044_), .A(_2415__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_3043_), );
  OAI21X1 OAI21X1_1258 (.Y(_3045_), .A(_3044_), .gnd(gnd), .vdd(vdd), .B(_3042_), .C(raddr1_2_bF_buf2_), );
  OAI21X1 OAI21X1_1259 (.Y(_3046_), .A(_1432_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf7_), .C(raddr1_1_bF_buf6_), );
  AOI21X1 AOI21X1_175 (.Y(_3047_), .A(regs_20__12_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf6_), .C(_3046_), );
  AND2X2 AND2X2_17 (.Y(_3048_), .A(regs_22__12_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf5_), );
  OAI21X1 OAI21X1_1260 (.Y(_3049_), .A(_1334_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf4_), .C(_2415__bF_buf0), );
  OAI21X1 OAI21X1_1261 (.Y(_3050_), .A(_3049_), .gnd(gnd), .vdd(vdd), .B(_3048_), .C(_2399__bF_buf1), );
  OAI22X1 OAI22X1_21 (.Y(_3051_), .A(_3041_), .gnd(gnd), .vdd(vdd), .B(_3045_), .C(_3050_), .D(_3047_), );
  INVX1 INVX1_65 (.Y(_3052_), .A(regs_29__12_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_457 (.Y(_3053_), .A(regs_28__12_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf3_), );
  OAI21X1 OAI21X1_1262 (.Y(_3054_), .A(_3052_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf2_), .C(_3053_), );
  MUX2X1 MUX2X1_118 (.Y(_3055_), .A(_3054_), .gnd(gnd), .vdd(vdd), .B(regs_30__12_), .S(raddr1_1_bF_buf5_), );
  NAND2X1 NAND2X1_458 (.Y(_3056_), .A(regs_26__12_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf1_), );
  OAI21X1 OAI21X1_1263 (.Y(_3057_), .A(_1167_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf0_), .C(_3056_), );
  INVX1 INVX1_66 (.Y(_3058_), .A(regs_25__12_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_459 (.Y(_3059_), .A(regs_24__12_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf96_), );
  OAI21X1 OAI21X1_1264 (.Y(_3060_), .A(_3058_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf95_), .C(_3059_), );
  MUX2X1 MUX2X1_119 (.Y(_3061_), .A(_3060_), .gnd(gnd), .vdd(vdd), .B(_3057_), .S(raddr1_1_bF_buf4_), );
  MUX2X1 MUX2X1_120 (.Y(_3062_), .A(_3061_), .gnd(gnd), .vdd(vdd), .B(_3055_), .S(raddr1_2_bF_buf1_), );
  MUX2X1 MUX2X1_121 (.Y(_3063_), .A(_3062_), .gnd(gnd), .vdd(vdd), .B(_3051_), .S(_2398__bF_buf1), );
  MUX2X1 MUX2X1_122 (.Y(_5511__12_), .A(_3039_), .gnd(gnd), .vdd(vdd), .B(_3063_), .S(raddr1_4_bF_buf2_), );
  INVX1 INVX1_67 (.Y(_3064_), .A(regs_5__13_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1265 (.Y(_3065_), .A(_3064_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf94_), .C(raddr1_1_bF_buf3_), );
  AOI21X1 AOI21X1_176 (.Y(_3066_), .A(regs_4__13_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf93_), .C(_3065_), );
  AND2X2 AND2X2_18 (.Y(_3067_), .A(regs_6__13_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf92_), );
  OAI21X1 OAI21X1_1266 (.Y(_3068_), .A(_2127_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf91_), .C(_2415__bF_buf8), );
  OAI21X1 OAI21X1_1267 (.Y(_3069_), .A(_3068_), .gnd(gnd), .vdd(vdd), .B(_3067_), .C(_2399__bF_buf0), );
  INVX1 INVX1_68 (.Y(_3070_), .A(regs_1__13_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1268 (.Y(_3071_), .A(_3070_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf90_), .C(raddr1_1_bF_buf2_), );
  AOI21X1 AOI21X1_177 (.Y(_3072_), .A(regs_0__13_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf89_), .C(_3071_), );
  INVX1 INVX1_69 (.Y(_3073_), .A(regs_3__13_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_164 (.Y(_3074_), .A(raddr1_0_bF_buf88_), .gnd(gnd), .vdd(vdd), .B(_3073_), );
  NAND2X1 NAND2X1_460 (.Y(_3075_), .A(regs_2__13_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf87_), );
  NAND2X1 NAND2X1_461 (.Y(_3076_), .A(_2415__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_3075_), );
  OAI21X1 OAI21X1_1269 (.Y(_3077_), .A(_3076_), .gnd(gnd), .vdd(vdd), .B(_3074_), .C(raddr1_2_bF_buf0_), );
  OAI22X1 OAI22X1_22 (.Y(_3078_), .A(_3072_), .gnd(gnd), .vdd(vdd), .B(_3077_), .C(_3069_), .D(_3066_), );
  NAND2X1 NAND2X1_462 (.Y(_3079_), .A(regs_10__13_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf86_), );
  OAI21X1 OAI21X1_1270 (.Y(_3080_), .A(_1928_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf85_), .C(_3079_), );
  NAND2X1 NAND2X1_463 (.Y(_3081_), .A(regs_8__13_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf84_), );
  OAI21X1 OAI21X1_1271 (.Y(_3082_), .A(_2026_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf83_), .C(_3081_), );
  MUX2X1 MUX2X1_123 (.Y(_3083_), .A(_3082_), .gnd(gnd), .vdd(vdd), .B(_3080_), .S(raddr1_1_bF_buf1_), );
  NAND2X1 NAND2X1_464 (.Y(_3084_), .A(regs_14__13_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf82_), );
  OAI21X1 OAI21X1_1272 (.Y(_3085_), .A(_1731_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf81_), .C(_3084_), );
  NAND2X1 NAND2X1_465 (.Y(_3086_), .A(regs_12__13_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf80_), );
  OAI21X1 OAI21X1_1273 (.Y(_3087_), .A(_1829_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf79_), .C(_3086_), );
  MUX2X1 MUX2X1_124 (.Y(_3088_), .A(_3087_), .gnd(gnd), .vdd(vdd), .B(_3085_), .S(raddr1_1_bF_buf0_), );
  MUX2X1 MUX2X1_125 (.Y(_3089_), .A(_3088_), .gnd(gnd), .vdd(vdd), .B(_3083_), .S(_2399__bF_buf8), );
  MUX2X1 MUX2X1_126 (.Y(_3090_), .A(_3089_), .gnd(gnd), .vdd(vdd), .B(_3078_), .S(_2398__bF_buf0), );
  OAI21X1 OAI21X1_1274 (.Y(_3091_), .A(_1631_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf78_), .C(raddr1_1_bF_buf14_bF_buf0_), );
  AOI21X1 AOI21X1_178 (.Y(_3092_), .A(regs_16__13_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf77_), .C(_3091_), );
  NOR2X1 NOR2X1_165 (.Y(_3093_), .A(raddr1_0_bF_buf76_), .gnd(gnd), .vdd(vdd), .B(_1533_), );
  NAND2X1 NAND2X1_466 (.Y(_3094_), .A(regs_18__13_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf75_), );
  NAND2X1 NAND2X1_467 (.Y(_3095_), .A(_2415__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_3094_), );
  OAI21X1 OAI21X1_1275 (.Y(_3096_), .A(_3095_), .gnd(gnd), .vdd(vdd), .B(_3093_), .C(raddr1_2_bF_buf10_), );
  OAI21X1 OAI21X1_1276 (.Y(_3097_), .A(_1434_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf74_), .C(raddr1_1_bF_buf13_bF_buf0_), );
  AOI21X1 AOI21X1_179 (.Y(_3098_), .A(regs_20__13_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf73_), .C(_3097_), );
  AND2X2 AND2X2_19 (.Y(_3099_), .A(regs_22__13_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf72_), );
  OAI21X1 OAI21X1_1277 (.Y(_3100_), .A(_1336_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf71_), .C(_2415__bF_buf5), );
  OAI21X1 OAI21X1_1278 (.Y(_3101_), .A(_3100_), .gnd(gnd), .vdd(vdd), .B(_3099_), .C(_2399__bF_buf7), );
  OAI22X1 OAI22X1_23 (.Y(_3102_), .A(_3092_), .gnd(gnd), .vdd(vdd), .B(_3096_), .C(_3101_), .D(_3098_), );
  INVX1 INVX1_70 (.Y(_3103_), .A(regs_29__13_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_468 (.Y(_3104_), .A(regs_28__13_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf70_), );
  OAI21X1 OAI21X1_1279 (.Y(_3105_), .A(_3103_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf69_), .C(_3104_), );
  MUX2X1 MUX2X1_127 (.Y(_3106_), .A(_3105_), .gnd(gnd), .vdd(vdd), .B(regs_30__13_), .S(raddr1_1_bF_buf12_bF_buf0_), );
  NAND2X1 NAND2X1_469 (.Y(_3107_), .A(regs_26__13_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf68_), );
  OAI21X1 OAI21X1_1280 (.Y(_3108_), .A(_1169_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf67_), .C(_3107_), );
  INVX1 INVX1_71 (.Y(_3109_), .A(regs_25__13_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_470 (.Y(_3110_), .A(regs_24__13_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf66_), );
  OAI21X1 OAI21X1_1281 (.Y(_3111_), .A(_3109_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf65_), .C(_3110_), );
  MUX2X1 MUX2X1_128 (.Y(_3112_), .A(_3111_), .gnd(gnd), .vdd(vdd), .B(_3108_), .S(raddr1_1_bF_buf11_bF_buf0_), );
  MUX2X1 MUX2X1_129 (.Y(_3113_), .A(_3112_), .gnd(gnd), .vdd(vdd), .B(_3106_), .S(raddr1_2_bF_buf9_), );
  MUX2X1 MUX2X1_130 (.Y(_3114_), .A(_3113_), .gnd(gnd), .vdd(vdd), .B(_3102_), .S(_2398__bF_buf7), );
  MUX2X1 MUX2X1_131 (.Y(_5511__13_), .A(_3090_), .gnd(gnd), .vdd(vdd), .B(_3114_), .S(raddr1_4_bF_buf1_), );
  NAND2X1 NAND2X1_471 (.Y(_3115_), .A(regs_22__14_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf64_), );
  OAI21X1 OAI21X1_1282 (.Y(_3116_), .A(_1338_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf63_), .C(_3115_), );
  NAND2X1 NAND2X1_472 (.Y(_3117_), .A(regs_20__14_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf62_), );
  OAI21X1 OAI21X1_1283 (.Y(_3118_), .A(_1436_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf61_), .C(_3117_), );
  MUX2X1 MUX2X1_132 (.Y(_3119_), .A(_3118_), .gnd(gnd), .vdd(vdd), .B(_3116_), .S(raddr1_1_bF_buf10_bF_buf0_), );
  NAND2X1 NAND2X1_473 (.Y(_3120_), .A(_2399__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_3119_), );
  NAND2X1 NAND2X1_474 (.Y(_3121_), .A(regs_18__14_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf60_), );
  OAI21X1 OAI21X1_1284 (.Y(_3122_), .A(_1535_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf59_), .C(_3121_), );
  NAND2X1 NAND2X1_475 (.Y(_3123_), .A(regs_16__14_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf58_), );
  OAI21X1 OAI21X1_1285 (.Y(_3124_), .A(_1633_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf57_), .C(_3123_), );
  MUX2X1 MUX2X1_133 (.Y(_3125_), .A(_3124_), .gnd(gnd), .vdd(vdd), .B(_3122_), .S(raddr1_1_bF_buf9_bF_buf0_), );
  AOI21X1 AOI21X1_180 (.Y(_3126_), .A(raddr1_2_bF_buf8_), .gnd(gnd), .vdd(vdd), .B(_3125_), .C(_2398__bF_buf6), );
  OAI21X1 OAI21X1_1286 (.Y(_3127_), .A(_1171_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf56_), .C(raddr1_2_bF_buf7_), );
  AOI21X1 AOI21X1_181 (.Y(_3128_), .A(regs_26__14_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf55_), .C(_3127_), );
  OAI21X1 OAI21X1_1287 (.Y(_3129_), .A(regs_30__14_), .gnd(gnd), .vdd(vdd), .B(raddr1_2_bF_buf6_), .C(_2415__bF_buf4), );
  INVX1 INVX1_72 (.Y(_3130_), .A(regs_25__14_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1288 (.Y(_3131_), .A(_3130_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf54_), .C(raddr1_2_bF_buf5_), );
  AOI21X1 AOI21X1_182 (.Y(_3132_), .A(regs_24__14_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf53_), .C(_3131_), );
  INVX1 INVX1_73 (.Y(_3133_), .A(regs_29__14_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_166 (.Y(_3134_), .A(raddr1_0_bF_buf52_), .gnd(gnd), .vdd(vdd), .B(_3133_), );
  NAND2X1 NAND2X1_476 (.Y(_3135_), .A(regs_28__14_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf51_), );
  NAND2X1 NAND2X1_477 (.Y(_3136_), .A(_2399__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_3135_), );
  OAI21X1 OAI21X1_1289 (.Y(_3137_), .A(_3136_), .gnd(gnd), .vdd(vdd), .B(_3134_), .C(raddr1_1_bF_buf8_), );
  OAI22X1 OAI22X1_24 (.Y(_3138_), .A(_3128_), .gnd(gnd), .vdd(vdd), .B(_3129_), .C(_3137_), .D(_3132_), );
  AOI22X1 AOI22X1_6 (.Y(_3139_), .A(_3138_), .gnd(gnd), .vdd(vdd), .B(_2398__bF_buf5), .C(_3120_), .D(_3126_), );
  INVX1 INVX1_74 (.Y(_3140_), .A(regs_5__14_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1290 (.Y(_3141_), .A(_3140_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf50_), .C(raddr1_1_bF_buf7_), );
  AOI21X1 AOI21X1_183 (.Y(_3142_), .A(regs_4__14_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf49_), .C(_3141_), );
  AND2X2 AND2X2_20 (.Y(_3143_), .A(regs_6__14_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf48_), );
  OAI21X1 OAI21X1_1291 (.Y(_3144_), .A(_2129_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf47_), .C(_2415__bF_buf3), );
  OAI21X1 OAI21X1_1292 (.Y(_3145_), .A(_3144_), .gnd(gnd), .vdd(vdd), .B(_3143_), .C(_2399__bF_buf4), );
  INVX1 INVX1_75 (.Y(_3146_), .A(regs_1__14_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1293 (.Y(_3147_), .A(_3146_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf46_), .C(raddr1_1_bF_buf6_), );
  AOI21X1 AOI21X1_184 (.Y(_3148_), .A(regs_0__14_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf45_), .C(_3147_), );
  INVX1 INVX1_76 (.Y(_3149_), .A(regs_3__14_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_167 (.Y(_3150_), .A(raddr1_0_bF_buf44_), .gnd(gnd), .vdd(vdd), .B(_3149_), );
  NAND2X1 NAND2X1_478 (.Y(_3151_), .A(regs_2__14_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf43_), );
  NAND2X1 NAND2X1_479 (.Y(_3152_), .A(_2415__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_3151_), );
  OAI21X1 OAI21X1_1294 (.Y(_3153_), .A(_3152_), .gnd(gnd), .vdd(vdd), .B(_3150_), .C(raddr1_2_bF_buf4_), );
  OAI22X1 OAI22X1_25 (.Y(_3154_), .A(_3148_), .gnd(gnd), .vdd(vdd), .B(_3153_), .C(_3145_), .D(_3142_), );
  NAND2X1 NAND2X1_480 (.Y(_3155_), .A(regs_10__14_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf42_), );
  OAI21X1 OAI21X1_1295 (.Y(_3156_), .A(_1930_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf41_), .C(_3155_), );
  NAND2X1 NAND2X1_481 (.Y(_3157_), .A(regs_8__14_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf40_), );
  OAI21X1 OAI21X1_1296 (.Y(_3158_), .A(_2028_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf39_), .C(_3157_), );
  MUX2X1 MUX2X1_134 (.Y(_3159_), .A(_3158_), .gnd(gnd), .vdd(vdd), .B(_3156_), .S(raddr1_1_bF_buf5_), );
  NAND2X1 NAND2X1_482 (.Y(_3160_), .A(regs_14__14_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf38_), );
  OAI21X1 OAI21X1_1297 (.Y(_3161_), .A(_1733_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf37_), .C(_3160_), );
  NAND2X1 NAND2X1_483 (.Y(_3162_), .A(regs_12__14_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf36_), );
  OAI21X1 OAI21X1_1298 (.Y(_3163_), .A(_1831_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf35_), .C(_3162_), );
  MUX2X1 MUX2X1_135 (.Y(_3164_), .A(_3163_), .gnd(gnd), .vdd(vdd), .B(_3161_), .S(raddr1_1_bF_buf4_), );
  MUX2X1 MUX2X1_136 (.Y(_3165_), .A(_3164_), .gnd(gnd), .vdd(vdd), .B(_3159_), .S(_2399__bF_buf3), );
  MUX2X1 MUX2X1_137 (.Y(_3166_), .A(_3165_), .gnd(gnd), .vdd(vdd), .B(_3154_), .S(_2398__bF_buf4), );
  MUX2X1 MUX2X1_138 (.Y(_5511__14_), .A(_3166_), .gnd(gnd), .vdd(vdd), .B(_3139_), .S(raddr1_4_bF_buf0_), );
  OAI21X1 OAI21X1_1299 (.Y(_3167_), .A(_1438_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf34_), .C(raddr1_1_bF_buf3_), );
  AOI21X1 AOI21X1_185 (.Y(_3168_), .A(regs_20__15_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf33_), .C(_3167_), );
  AND2X2 AND2X2_21 (.Y(_3169_), .A(regs_22__15_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf32_), );
  OAI21X1 OAI21X1_1300 (.Y(_3170_), .A(_1340_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf31_), .C(_2415__bF_buf1), );
  OAI21X1 OAI21X1_1301 (.Y(_3171_), .A(_3170_), .gnd(gnd), .vdd(vdd), .B(_3169_), .C(_2399__bF_buf2), );
  OAI21X1 OAI21X1_1302 (.Y(_3172_), .A(_1635_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf30_), .C(raddr1_1_bF_buf2_), );
  AOI21X1 AOI21X1_186 (.Y(_3173_), .A(regs_16__15_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf29_), .C(_3172_), );
  NOR2X1 NOR2X1_168 (.Y(_3174_), .A(raddr1_0_bF_buf28_), .gnd(gnd), .vdd(vdd), .B(_1537_), );
  NAND2X1 NAND2X1_484 (.Y(_3175_), .A(regs_18__15_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf27_), );
  NAND2X1 NAND2X1_485 (.Y(_3176_), .A(_2415__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_3175_), );
  OAI21X1 OAI21X1_1303 (.Y(_3177_), .A(_3176_), .gnd(gnd), .vdd(vdd), .B(_3174_), .C(raddr1_2_bF_buf3_), );
  OAI22X1 OAI22X1_26 (.Y(_3178_), .A(_3173_), .gnd(gnd), .vdd(vdd), .B(_3177_), .C(_3171_), .D(_3168_), );
  INVX1 INVX1_77 (.Y(_3179_), .A(regs_29__15_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_486 (.Y(_3180_), .A(regs_28__15_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf26_), );
  OAI21X1 OAI21X1_1304 (.Y(_3181_), .A(_3179_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf25_), .C(_3180_), );
  MUX2X1 MUX2X1_139 (.Y(_3182_), .A(_3181_), .gnd(gnd), .vdd(vdd), .B(regs_30__15_), .S(raddr1_1_bF_buf1_), );
  NAND2X1 NAND2X1_487 (.Y(_3183_), .A(regs_26__15_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf24_), );
  OAI21X1 OAI21X1_1305 (.Y(_3184_), .A(_1173_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf23_), .C(_3183_), );
  INVX1 INVX1_78 (.Y(_3185_), .A(regs_25__15_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_488 (.Y(_3186_), .A(regs_24__15_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf22_), );
  OAI21X1 OAI21X1_1306 (.Y(_3187_), .A(_3185_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf21_), .C(_3186_), );
  MUX2X1 MUX2X1_140 (.Y(_3188_), .A(_3187_), .gnd(gnd), .vdd(vdd), .B(_3184_), .S(raddr1_1_bF_buf0_), );
  MUX2X1 MUX2X1_141 (.Y(_3189_), .A(_3188_), .gnd(gnd), .vdd(vdd), .B(_3182_), .S(raddr1_2_bF_buf2_), );
  MUX2X1 MUX2X1_142 (.Y(_3190_), .A(_3189_), .gnd(gnd), .vdd(vdd), .B(_3178_), .S(_2398__bF_buf3), );
  NAND2X1 NAND2X1_489 (.Y(_3191_), .A(regs_6__15_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf20_), );
  OAI21X1 OAI21X1_1307 (.Y(_3192_), .A(_2131_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf19_), .C(_3191_), );
  INVX1 INVX1_79 (.Y(_3193_), .A(regs_5__15_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_490 (.Y(_3194_), .A(regs_4__15_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf18_), );
  OAI21X1 OAI21X1_1308 (.Y(_3195_), .A(_3193_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf17_), .C(_3194_), );
  MUX2X1 MUX2X1_143 (.Y(_3196_), .A(_3195_), .gnd(gnd), .vdd(vdd), .B(_3192_), .S(raddr1_1_bF_buf14_bF_buf3_), );
  INVX1 INVX1_80 (.Y(_3197_), .A(regs_3__15_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_491 (.Y(_3198_), .A(regs_2__15_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf16_), );
  OAI21X1 OAI21X1_1309 (.Y(_3199_), .A(_3197_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf15_), .C(_3198_), );
  INVX1 INVX1_81 (.Y(_3200_), .A(regs_1__15_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_492 (.Y(_3201_), .A(regs_0__15_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf14_), );
  OAI21X1 OAI21X1_1310 (.Y(_3202_), .A(_3200_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf13_), .C(_3201_), );
  MUX2X1 MUX2X1_144 (.Y(_3203_), .A(_3202_), .gnd(gnd), .vdd(vdd), .B(_3199_), .S(raddr1_1_bF_buf13_bF_buf3_), );
  MUX2X1 MUX2X1_145 (.Y(_3204_), .A(_3203_), .gnd(gnd), .vdd(vdd), .B(_3196_), .S(raddr1_2_bF_buf1_), );
  NAND2X1 NAND2X1_493 (.Y(_3205_), .A(regs_14__15_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf12_), );
  OAI21X1 OAI21X1_1311 (.Y(_3206_), .A(_1735_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf11_), .C(_3205_), );
  NAND2X1 NAND2X1_494 (.Y(_3207_), .A(regs_12__15_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf10_), );
  OAI21X1 OAI21X1_1312 (.Y(_3208_), .A(_1833_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf9_), .C(_3207_), );
  MUX2X1 MUX2X1_146 (.Y(_3209_), .A(_3208_), .gnd(gnd), .vdd(vdd), .B(_3206_), .S(raddr1_1_bF_buf12_bF_buf3_), );
  NAND2X1 NAND2X1_495 (.Y(_3210_), .A(regs_10__15_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf8_), );
  OAI21X1 OAI21X1_1313 (.Y(_3211_), .A(_1932_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf7_), .C(_3210_), );
  NAND2X1 NAND2X1_496 (.Y(_3212_), .A(regs_8__15_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf6_), );
  OAI21X1 OAI21X1_1314 (.Y(_3213_), .A(_2030_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf5_), .C(_3212_), );
  MUX2X1 MUX2X1_147 (.Y(_3214_), .A(_3213_), .gnd(gnd), .vdd(vdd), .B(_3211_), .S(raddr1_1_bF_buf11_bF_buf3_), );
  MUX2X1 MUX2X1_148 (.Y(_3215_), .A(_3214_), .gnd(gnd), .vdd(vdd), .B(_3209_), .S(raddr1_2_bF_buf0_), );
  MUX2X1 MUX2X1_149 (.Y(_3216_), .A(_3215_), .gnd(gnd), .vdd(vdd), .B(_3204_), .S(_2398__bF_buf2), );
  MUX2X1 MUX2X1_150 (.Y(_5511__15_), .A(_3216_), .gnd(gnd), .vdd(vdd), .B(_3190_), .S(raddr1_4_bF_buf4_), );
  NAND2X1 NAND2X1_497 (.Y(_3217_), .A(regs_22__16_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf4_), );
  OAI21X1 OAI21X1_1315 (.Y(_3218_), .A(_1342_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf3_), .C(_3217_), );
  NAND2X1 NAND2X1_498 (.Y(_3219_), .A(regs_20__16_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf2_), );
  OAI21X1 OAI21X1_1316 (.Y(_3220_), .A(_1440_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf1_), .C(_3219_), );
  MUX2X1 MUX2X1_151 (.Y(_3221_), .A(_3220_), .gnd(gnd), .vdd(vdd), .B(_3218_), .S(raddr1_1_bF_buf10_bF_buf3_), );
  NAND2X1 NAND2X1_499 (.Y(_3222_), .A(_2399__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_3221_), );
  NAND2X1 NAND2X1_500 (.Y(_3223_), .A(regs_18__16_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf0_), );
  OAI21X1 OAI21X1_1317 (.Y(_3224_), .A(_1539_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf96_), .C(_3223_), );
  NAND2X1 NAND2X1_501 (.Y(_3225_), .A(regs_16__16_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf95_), );
  OAI21X1 OAI21X1_1318 (.Y(_3226_), .A(_1637_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf94_), .C(_3225_), );
  MUX2X1 MUX2X1_152 (.Y(_3227_), .A(_3226_), .gnd(gnd), .vdd(vdd), .B(_3224_), .S(raddr1_1_bF_buf9_bF_buf3_), );
  AOI21X1 AOI21X1_187 (.Y(_3228_), .A(raddr1_2_bF_buf10_), .gnd(gnd), .vdd(vdd), .B(_3227_), .C(_2398__bF_buf1), );
  OAI21X1 OAI21X1_1319 (.Y(_3229_), .A(_1175_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf93_), .C(raddr1_2_bF_buf9_), );
  AOI21X1 AOI21X1_188 (.Y(_3230_), .A(regs_26__16_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf92_), .C(_3229_), );
  OAI21X1 OAI21X1_1320 (.Y(_3231_), .A(regs_30__16_), .gnd(gnd), .vdd(vdd), .B(raddr1_2_bF_buf8_), .C(_2415__bF_buf8), );
  INVX1 INVX1_82 (.Y(_3232_), .A(regs_25__16_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1321 (.Y(_3233_), .A(_3232_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf91_), .C(raddr1_2_bF_buf7_), );
  AOI21X1 AOI21X1_189 (.Y(_3234_), .A(regs_24__16_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf90_), .C(_3233_), );
  INVX1 INVX1_83 (.Y(_3235_), .A(regs_29__16_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_169 (.Y(_3236_), .A(raddr1_0_bF_buf89_), .gnd(gnd), .vdd(vdd), .B(_3235_), );
  NAND2X1 NAND2X1_502 (.Y(_3237_), .A(regs_28__16_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf88_), );
  NAND2X1 NAND2X1_503 (.Y(_3238_), .A(_2399__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_3237_), );
  OAI21X1 OAI21X1_1322 (.Y(_3239_), .A(_3238_), .gnd(gnd), .vdd(vdd), .B(_3236_), .C(raddr1_1_bF_buf8_), );
  OAI22X1 OAI22X1_27 (.Y(_3240_), .A(_3230_), .gnd(gnd), .vdd(vdd), .B(_3231_), .C(_3239_), .D(_3234_), );
  AOI22X1 AOI22X1_7 (.Y(_3241_), .A(_3240_), .gnd(gnd), .vdd(vdd), .B(_2398__bF_buf0), .C(_3222_), .D(_3228_), );
  INVX1 INVX1_84 (.Y(_3242_), .A(regs_5__16_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1323 (.Y(_3243_), .A(_3242_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf87_), .C(raddr1_1_bF_buf7_), );
  AOI21X1 AOI21X1_190 (.Y(_3244_), .A(regs_4__16_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf86_), .C(_3243_), );
  AND2X2 AND2X2_22 (.Y(_3245_), .A(regs_6__16_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf85_), );
  OAI21X1 OAI21X1_1324 (.Y(_3246_), .A(_2133_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf84_), .C(_2415__bF_buf7), );
  OAI21X1 OAI21X1_1325 (.Y(_3247_), .A(_3246_), .gnd(gnd), .vdd(vdd), .B(_3245_), .C(_2399__bF_buf8), );
  INVX1 INVX1_85 (.Y(_3248_), .A(regs_1__16_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1326 (.Y(_3249_), .A(_3248_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf83_), .C(raddr1_1_bF_buf6_), );
  AOI21X1 AOI21X1_191 (.Y(_3250_), .A(regs_0__16_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf82_), .C(_3249_), );
  INVX1 INVX1_86 (.Y(_3251_), .A(regs_3__16_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_170 (.Y(_3252_), .A(raddr1_0_bF_buf81_), .gnd(gnd), .vdd(vdd), .B(_3251_), );
  NAND2X1 NAND2X1_504 (.Y(_3253_), .A(regs_2__16_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf80_), );
  NAND2X1 NAND2X1_505 (.Y(_3254_), .A(_2415__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_3253_), );
  OAI21X1 OAI21X1_1327 (.Y(_3255_), .A(_3254_), .gnd(gnd), .vdd(vdd), .B(_3252_), .C(raddr1_2_bF_buf6_), );
  OAI22X1 OAI22X1_28 (.Y(_3256_), .A(_3250_), .gnd(gnd), .vdd(vdd), .B(_3255_), .C(_3247_), .D(_3244_), );
  NAND2X1 NAND2X1_506 (.Y(_3257_), .A(regs_10__16_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf79_), );
  OAI21X1 OAI21X1_1328 (.Y(_3258_), .A(_1934_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf78_), .C(_3257_), );
  NAND2X1 NAND2X1_507 (.Y(_3259_), .A(regs_8__16_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf77_), );
  OAI21X1 OAI21X1_1329 (.Y(_3260_), .A(_2032_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf76_), .C(_3259_), );
  MUX2X1 MUX2X1_153 (.Y(_3261_), .A(_3260_), .gnd(gnd), .vdd(vdd), .B(_3258_), .S(raddr1_1_bF_buf5_), );
  NAND2X1 NAND2X1_508 (.Y(_3262_), .A(regs_14__16_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf75_), );
  OAI21X1 OAI21X1_1330 (.Y(_3263_), .A(_1737_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf74_), .C(_3262_), );
  NAND2X1 NAND2X1_509 (.Y(_3264_), .A(regs_12__16_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf73_), );
  OAI21X1 OAI21X1_1331 (.Y(_3265_), .A(_1835_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf72_), .C(_3264_), );
  MUX2X1 MUX2X1_154 (.Y(_3266_), .A(_3265_), .gnd(gnd), .vdd(vdd), .B(_3263_), .S(raddr1_1_bF_buf4_), );
  MUX2X1 MUX2X1_155 (.Y(_3267_), .A(_3266_), .gnd(gnd), .vdd(vdd), .B(_3261_), .S(_2399__bF_buf7), );
  MUX2X1 MUX2X1_156 (.Y(_3268_), .A(_3267_), .gnd(gnd), .vdd(vdd), .B(_3256_), .S(_2398__bF_buf7), );
  MUX2X1 MUX2X1_157 (.Y(_5511__16_), .A(_3268_), .gnd(gnd), .vdd(vdd), .B(_3241_), .S(raddr1_4_bF_buf3_), );
  NAND2X1 NAND2X1_510 (.Y(_3269_), .A(regs_22__17_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf71_), );
  OAI21X1 OAI21X1_1332 (.Y(_3270_), .A(_1344_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf70_), .C(_3269_), );
  NAND2X1 NAND2X1_511 (.Y(_3271_), .A(regs_20__17_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf69_), );
  OAI21X1 OAI21X1_1333 (.Y(_3272_), .A(_1442_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf68_), .C(_3271_), );
  MUX2X1 MUX2X1_158 (.Y(_3273_), .A(_3272_), .gnd(gnd), .vdd(vdd), .B(_3270_), .S(raddr1_1_bF_buf3_), );
  NAND2X1 NAND2X1_512 (.Y(_3274_), .A(_2399__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_3273_), );
  NAND2X1 NAND2X1_513 (.Y(_3275_), .A(regs_18__17_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf67_), );
  OAI21X1 OAI21X1_1334 (.Y(_3276_), .A(_1541_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf66_), .C(_3275_), );
  NAND2X1 NAND2X1_514 (.Y(_3277_), .A(regs_16__17_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf65_), );
  OAI21X1 OAI21X1_1335 (.Y(_3278_), .A(_1639_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf64_), .C(_3277_), );
  MUX2X1 MUX2X1_159 (.Y(_3279_), .A(_3278_), .gnd(gnd), .vdd(vdd), .B(_3276_), .S(raddr1_1_bF_buf2_), );
  AOI21X1 AOI21X1_192 (.Y(_3280_), .A(raddr1_2_bF_buf5_), .gnd(gnd), .vdd(vdd), .B(_3279_), .C(_2398__bF_buf6), );
  OAI21X1 OAI21X1_1336 (.Y(_3281_), .A(_1177_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf63_), .C(raddr1_2_bF_buf4_), );
  AOI21X1 AOI21X1_193 (.Y(_3282_), .A(regs_26__17_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf62_), .C(_3281_), );
  OAI21X1 OAI21X1_1337 (.Y(_3283_), .A(regs_30__17_), .gnd(gnd), .vdd(vdd), .B(raddr1_2_bF_buf3_), .C(_2415__bF_buf5), );
  INVX1 INVX1_87 (.Y(_3284_), .A(regs_25__17_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1338 (.Y(_3285_), .A(_3284_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf61_), .C(raddr1_2_bF_buf2_), );
  AOI21X1 AOI21X1_194 (.Y(_3286_), .A(regs_24__17_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf60_), .C(_3285_), );
  INVX1 INVX1_88 (.Y(_3287_), .A(regs_29__17_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_171 (.Y(_3288_), .A(raddr1_0_bF_buf59_), .gnd(gnd), .vdd(vdd), .B(_3287_), );
  NAND2X1 NAND2X1_515 (.Y(_3289_), .A(regs_28__17_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf58_), );
  NAND2X1 NAND2X1_516 (.Y(_3290_), .A(_2399__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_3289_), );
  OAI21X1 OAI21X1_1339 (.Y(_3291_), .A(_3290_), .gnd(gnd), .vdd(vdd), .B(_3288_), .C(raddr1_1_bF_buf1_), );
  OAI22X1 OAI22X1_29 (.Y(_3292_), .A(_3282_), .gnd(gnd), .vdd(vdd), .B(_3283_), .C(_3291_), .D(_3286_), );
  AOI22X1 AOI22X1_8 (.Y(_3293_), .A(_3292_), .gnd(gnd), .vdd(vdd), .B(_2398__bF_buf5), .C(_3274_), .D(_3280_), );
  INVX1 INVX1_89 (.Y(_3294_), .A(regs_5__17_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1340 (.Y(_3295_), .A(_3294_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf57_), .C(raddr1_1_bF_buf0_), );
  AOI21X1 AOI21X1_195 (.Y(_3296_), .A(regs_4__17_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf56_), .C(_3295_), );
  AND2X2 AND2X2_23 (.Y(_3297_), .A(regs_6__17_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf55_), );
  OAI21X1 OAI21X1_1341 (.Y(_3298_), .A(_2135_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf54_), .C(_2415__bF_buf4), );
  OAI21X1 OAI21X1_1342 (.Y(_3299_), .A(_3298_), .gnd(gnd), .vdd(vdd), .B(_3297_), .C(_2399__bF_buf4), );
  INVX1 INVX1_90 (.Y(_3300_), .A(regs_1__17_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1343 (.Y(_3301_), .A(_3300_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf53_), .C(raddr1_1_bF_buf14_bF_buf2_), );
  AOI21X1 AOI21X1_196 (.Y(_3302_), .A(regs_0__17_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf52_), .C(_3301_), );
  INVX1 INVX1_91 (.Y(_3303_), .A(regs_3__17_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_172 (.Y(_3304_), .A(raddr1_0_bF_buf51_), .gnd(gnd), .vdd(vdd), .B(_3303_), );
  NAND2X1 NAND2X1_517 (.Y(_3305_), .A(regs_2__17_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf50_), );
  NAND2X1 NAND2X1_518 (.Y(_3306_), .A(_2415__bF_buf3), .gnd(gnd), .vdd(vdd), .B(_3305_), );
  OAI21X1 OAI21X1_1344 (.Y(_3307_), .A(_3306_), .gnd(gnd), .vdd(vdd), .B(_3304_), .C(raddr1_2_bF_buf1_), );
  OAI22X1 OAI22X1_30 (.Y(_3308_), .A(_3302_), .gnd(gnd), .vdd(vdd), .B(_3307_), .C(_3299_), .D(_3296_), );
  NAND2X1 NAND2X1_519 (.Y(_3309_), .A(regs_10__17_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf49_), );
  OAI21X1 OAI21X1_1345 (.Y(_3310_), .A(_1936_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf48_), .C(_3309_), );
  NAND2X1 NAND2X1_520 (.Y(_3311_), .A(regs_8__17_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf47_), );
  OAI21X1 OAI21X1_1346 (.Y(_3312_), .A(_2034_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf46_), .C(_3311_), );
  MUX2X1 MUX2X1_160 (.Y(_3313_), .A(_3312_), .gnd(gnd), .vdd(vdd), .B(_3310_), .S(raddr1_1_bF_buf13_bF_buf2_), );
  NAND2X1 NAND2X1_521 (.Y(_3314_), .A(regs_14__17_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf45_), );
  OAI21X1 OAI21X1_1347 (.Y(_3315_), .A(_1739_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf44_), .C(_3314_), );
  NAND2X1 NAND2X1_522 (.Y(_3316_), .A(regs_12__17_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf43_), );
  OAI21X1 OAI21X1_1348 (.Y(_3317_), .A(_1837_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf42_), .C(_3316_), );
  MUX2X1 MUX2X1_161 (.Y(_3318_), .A(_3317_), .gnd(gnd), .vdd(vdd), .B(_3315_), .S(raddr1_1_bF_buf12_bF_buf2_), );
  MUX2X1 MUX2X1_162 (.Y(_3319_), .A(_3318_), .gnd(gnd), .vdd(vdd), .B(_3313_), .S(_2399__bF_buf3), );
  MUX2X1 MUX2X1_163 (.Y(_3320_), .A(_3319_), .gnd(gnd), .vdd(vdd), .B(_3308_), .S(_2398__bF_buf4), );
  MUX2X1 MUX2X1_164 (.Y(_5511__17_), .A(_3320_), .gnd(gnd), .vdd(vdd), .B(_3293_), .S(raddr1_4_bF_buf2_), );
  INVX1 INVX1_92 (.Y(_3321_), .A(regs_5__18_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1349 (.Y(_3322_), .A(_3321_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf41_), .C(raddr1_1_bF_buf11_bF_buf2_), );
  AOI21X1 AOI21X1_197 (.Y(_3323_), .A(regs_4__18_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf40_), .C(_3322_), );
  AND2X2 AND2X2_24 (.Y(_3324_), .A(regs_6__18_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf39_), );
  OAI21X1 OAI21X1_1350 (.Y(_3325_), .A(_2137_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf38_), .C(_2415__bF_buf2), );
  OAI21X1 OAI21X1_1351 (.Y(_3326_), .A(_3325_), .gnd(gnd), .vdd(vdd), .B(_3324_), .C(_2399__bF_buf2), );
  INVX1 INVX1_93 (.Y(_3327_), .A(regs_1__18_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1352 (.Y(_3328_), .A(_3327_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf37_), .C(raddr1_1_bF_buf10_bF_buf2_), );
  AOI21X1 AOI21X1_198 (.Y(_3329_), .A(regs_0__18_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf36_), .C(_3328_), );
  INVX1 INVX1_94 (.Y(_3330_), .A(regs_3__18_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_173 (.Y(_3331_), .A(raddr1_0_bF_buf35_), .gnd(gnd), .vdd(vdd), .B(_3330_), );
  NAND2X1 NAND2X1_523 (.Y(_3332_), .A(regs_2__18_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf34_), );
  NAND2X1 NAND2X1_524 (.Y(_3333_), .A(_2415__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_3332_), );
  OAI21X1 OAI21X1_1353 (.Y(_3334_), .A(_3333_), .gnd(gnd), .vdd(vdd), .B(_3331_), .C(raddr1_2_bF_buf0_), );
  OAI22X1 OAI22X1_31 (.Y(_3335_), .A(_3329_), .gnd(gnd), .vdd(vdd), .B(_3334_), .C(_3326_), .D(_3323_), );
  NAND2X1 NAND2X1_525 (.Y(_3336_), .A(regs_10__18_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf33_), );
  OAI21X1 OAI21X1_1354 (.Y(_3337_), .A(_1938_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf32_), .C(_3336_), );
  NAND2X1 NAND2X1_526 (.Y(_3338_), .A(regs_8__18_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf31_), );
  OAI21X1 OAI21X1_1355 (.Y(_3339_), .A(_2036_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf30_), .C(_3338_), );
  MUX2X1 MUX2X1_165 (.Y(_3340_), .A(_3339_), .gnd(gnd), .vdd(vdd), .B(_3337_), .S(raddr1_1_bF_buf9_bF_buf2_), );
  NAND2X1 NAND2X1_527 (.Y(_3341_), .A(regs_14__18_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf29_), );
  OAI21X1 OAI21X1_1356 (.Y(_3342_), .A(_1741_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf28_), .C(_3341_), );
  NAND2X1 NAND2X1_528 (.Y(_3343_), .A(regs_12__18_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf27_), );
  OAI21X1 OAI21X1_1357 (.Y(_3344_), .A(_1839_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf26_), .C(_3343_), );
  MUX2X1 MUX2X1_166 (.Y(_3345_), .A(_3344_), .gnd(gnd), .vdd(vdd), .B(_3342_), .S(raddr1_1_bF_buf8_), );
  MUX2X1 MUX2X1_167 (.Y(_3346_), .A(_3345_), .gnd(gnd), .vdd(vdd), .B(_3340_), .S(_2399__bF_buf1), );
  MUX2X1 MUX2X1_168 (.Y(_3347_), .A(_3346_), .gnd(gnd), .vdd(vdd), .B(_3335_), .S(_2398__bF_buf3), );
  OAI21X1 OAI21X1_1358 (.Y(_3348_), .A(_1641_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf25_), .C(raddr1_1_bF_buf7_), );
  AOI21X1 AOI21X1_199 (.Y(_3349_), .A(regs_16__18_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf24_), .C(_3348_), );
  NOR2X1 NOR2X1_174 (.Y(_3350_), .A(raddr1_0_bF_buf23_), .gnd(gnd), .vdd(vdd), .B(_1543_), );
  NAND2X1 NAND2X1_529 (.Y(_3351_), .A(regs_18__18_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf22_), );
  NAND2X1 NAND2X1_530 (.Y(_3352_), .A(_2415__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_3351_), );
  OAI21X1 OAI21X1_1359 (.Y(_3353_), .A(_3352_), .gnd(gnd), .vdd(vdd), .B(_3350_), .C(raddr1_2_bF_buf10_), );
  OAI21X1 OAI21X1_1360 (.Y(_3354_), .A(_1444_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf21_), .C(raddr1_1_bF_buf6_), );
  AOI21X1 AOI21X1_200 (.Y(_3355_), .A(regs_20__18_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf20_), .C(_3354_), );
  AND2X2 AND2X2_25 (.Y(_3356_), .A(regs_22__18_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf19_), );
  OAI21X1 OAI21X1_1361 (.Y(_3357_), .A(_1346_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf18_), .C(_2415__bF_buf8), );
  OAI21X1 OAI21X1_1362 (.Y(_3358_), .A(_3357_), .gnd(gnd), .vdd(vdd), .B(_3356_), .C(_2399__bF_buf0), );
  OAI22X1 OAI22X1_32 (.Y(_3359_), .A(_3349_), .gnd(gnd), .vdd(vdd), .B(_3353_), .C(_3358_), .D(_3355_), );
  INVX1 INVX1_95 (.Y(_3360_), .A(regs_29__18_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_531 (.Y(_3361_), .A(regs_28__18_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf17_), );
  OAI21X1 OAI21X1_1363 (.Y(_3362_), .A(_3360_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf16_), .C(_3361_), );
  MUX2X1 MUX2X1_169 (.Y(_3363_), .A(_3362_), .gnd(gnd), .vdd(vdd), .B(regs_30__18_), .S(raddr1_1_bF_buf5_), );
  NAND2X1 NAND2X1_532 (.Y(_3364_), .A(regs_26__18_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf15_), );
  OAI21X1 OAI21X1_1364 (.Y(_3365_), .A(_1179_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf14_), .C(_3364_), );
  INVX1 INVX1_96 (.Y(_3366_), .A(regs_25__18_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_533 (.Y(_3367_), .A(regs_24__18_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf13_), );
  OAI21X1 OAI21X1_1365 (.Y(_3368_), .A(_3366_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf12_), .C(_3367_), );
  MUX2X1 MUX2X1_170 (.Y(_3369_), .A(_3368_), .gnd(gnd), .vdd(vdd), .B(_3365_), .S(raddr1_1_bF_buf4_), );
  MUX2X1 MUX2X1_171 (.Y(_3370_), .A(_3369_), .gnd(gnd), .vdd(vdd), .B(_3363_), .S(raddr1_2_bF_buf9_), );
  MUX2X1 MUX2X1_172 (.Y(_3371_), .A(_3370_), .gnd(gnd), .vdd(vdd), .B(_3359_), .S(_2398__bF_buf2), );
  MUX2X1 MUX2X1_173 (.Y(_5511__18_), .A(_3347_), .gnd(gnd), .vdd(vdd), .B(_3371_), .S(raddr1_4_bF_buf1_), );
  NAND2X1 NAND2X1_534 (.Y(_3372_), .A(regs_22__19_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf11_), );
  OAI21X1 OAI21X1_1366 (.Y(_3373_), .A(_1348_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf10_), .C(_3372_), );
  NAND2X1 NAND2X1_535 (.Y(_3374_), .A(regs_20__19_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf9_), );
  OAI21X1 OAI21X1_1367 (.Y(_3375_), .A(_1446_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf8_), .C(_3374_), );
  MUX2X1 MUX2X1_174 (.Y(_3376_), .A(_3375_), .gnd(gnd), .vdd(vdd), .B(_3373_), .S(raddr1_1_bF_buf3_), );
  NAND2X1 NAND2X1_536 (.Y(_3377_), .A(_2399__bF_buf8), .gnd(gnd), .vdd(vdd), .B(_3376_), );
  NAND2X1 NAND2X1_537 (.Y(_3378_), .A(regs_18__19_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf7_), );
  OAI21X1 OAI21X1_1368 (.Y(_3379_), .A(_1545_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf6_), .C(_3378_), );
  NAND2X1 NAND2X1_538 (.Y(_3380_), .A(regs_16__19_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf5_), );
  OAI21X1 OAI21X1_1369 (.Y(_3381_), .A(_1643_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf4_), .C(_3380_), );
  MUX2X1 MUX2X1_175 (.Y(_3382_), .A(_3381_), .gnd(gnd), .vdd(vdd), .B(_3379_), .S(raddr1_1_bF_buf2_), );
  AOI21X1 AOI21X1_201 (.Y(_3383_), .A(raddr1_2_bF_buf8_), .gnd(gnd), .vdd(vdd), .B(_3382_), .C(_2398__bF_buf1), );
  OAI21X1 OAI21X1_1370 (.Y(_3384_), .A(_1181_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf3_), .C(raddr1_2_bF_buf7_), );
  AOI21X1 AOI21X1_202 (.Y(_3385_), .A(regs_26__19_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf2_), .C(_3384_), );
  OAI21X1 OAI21X1_1371 (.Y(_3386_), .A(regs_30__19_), .gnd(gnd), .vdd(vdd), .B(raddr1_2_bF_buf6_), .C(_2415__bF_buf7), );
  INVX1 INVX1_97 (.Y(_3387_), .A(regs_25__19_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1372 (.Y(_3388_), .A(_3387_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf1_), .C(raddr1_2_bF_buf5_), );
  AOI21X1 AOI21X1_203 (.Y(_3389_), .A(regs_24__19_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf0_), .C(_3388_), );
  INVX1 INVX1_98 (.Y(_3390_), .A(regs_29__19_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_175 (.Y(_3391_), .A(raddr1_0_bF_buf96_), .gnd(gnd), .vdd(vdd), .B(_3390_), );
  NAND2X1 NAND2X1_539 (.Y(_3392_), .A(regs_28__19_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf95_), );
  NAND2X1 NAND2X1_540 (.Y(_3393_), .A(_2399__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_3392_), );
  OAI21X1 OAI21X1_1373 (.Y(_3394_), .A(_3393_), .gnd(gnd), .vdd(vdd), .B(_3391_), .C(raddr1_1_bF_buf1_), );
  OAI22X1 OAI22X1_33 (.Y(_3395_), .A(_3385_), .gnd(gnd), .vdd(vdd), .B(_3386_), .C(_3394_), .D(_3389_), );
  AOI22X1 AOI22X1_9 (.Y(_3396_), .A(_3395_), .gnd(gnd), .vdd(vdd), .B(_2398__bF_buf0), .C(_3377_), .D(_3383_), );
  NAND2X1 NAND2X1_541 (.Y(_3397_), .A(regs_6__19_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf94_), );
  OAI21X1 OAI21X1_1374 (.Y(_3398_), .A(_2139_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf93_), .C(_3397_), );
  INVX1 INVX1_99 (.Y(_3399_), .A(regs_5__19_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_542 (.Y(_3400_), .A(regs_4__19_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf92_), );
  OAI21X1 OAI21X1_1375 (.Y(_3401_), .A(_3399_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf91_), .C(_3400_), );
  MUX2X1 MUX2X1_176 (.Y(_3402_), .A(_3401_), .gnd(gnd), .vdd(vdd), .B(_3398_), .S(raddr1_1_bF_buf0_), );
  INVX1 INVX1_100 (.Y(_3403_), .A(regs_3__19_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_543 (.Y(_3404_), .A(regs_2__19_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf90_), );
  OAI21X1 OAI21X1_1376 (.Y(_3405_), .A(_3403_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf89_), .C(_3404_), );
  INVX1 INVX1_101 (.Y(_3406_), .A(regs_1__19_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_544 (.Y(_3407_), .A(regs_0__19_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf88_), );
  OAI21X1 OAI21X1_1377 (.Y(_3408_), .A(_3406_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf87_), .C(_3407_), );
  MUX2X1 MUX2X1_177 (.Y(_3409_), .A(_3408_), .gnd(gnd), .vdd(vdd), .B(_3405_), .S(raddr1_1_bF_buf14_bF_buf1_), );
  MUX2X1 MUX2X1_178 (.Y(_3410_), .A(_3409_), .gnd(gnd), .vdd(vdd), .B(_3402_), .S(raddr1_2_bF_buf4_), );
  NAND2X1 NAND2X1_545 (.Y(_3411_), .A(regs_10__19_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf86_), );
  OAI21X1 OAI21X1_1378 (.Y(_3412_), .A(_1940_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf85_), .C(_3411_), );
  NAND2X1 NAND2X1_546 (.Y(_3413_), .A(regs_8__19_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf84_), );
  OAI21X1 OAI21X1_1379 (.Y(_3414_), .A(_2038_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf83_), .C(_3413_), );
  MUX2X1 MUX2X1_179 (.Y(_3415_), .A(_3414_), .gnd(gnd), .vdd(vdd), .B(_3412_), .S(raddr1_1_bF_buf13_bF_buf1_), );
  NAND2X1 NAND2X1_547 (.Y(_3416_), .A(regs_14__19_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf82_), );
  OAI21X1 OAI21X1_1380 (.Y(_3417_), .A(_1743_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf81_), .C(_3416_), );
  NAND2X1 NAND2X1_548 (.Y(_3418_), .A(regs_12__19_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf80_), );
  OAI21X1 OAI21X1_1381 (.Y(_3419_), .A(_1841_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf79_), .C(_3418_), );
  MUX2X1 MUX2X1_180 (.Y(_3420_), .A(_3419_), .gnd(gnd), .vdd(vdd), .B(_3417_), .S(raddr1_1_bF_buf12_bF_buf1_), );
  MUX2X1 MUX2X1_181 (.Y(_3421_), .A(_3420_), .gnd(gnd), .vdd(vdd), .B(_3415_), .S(_2399__bF_buf6), );
  MUX2X1 MUX2X1_182 (.Y(_3422_), .A(_3421_), .gnd(gnd), .vdd(vdd), .B(_3410_), .S(_2398__bF_buf7), );
  MUX2X1 MUX2X1_183 (.Y(_5511__19_), .A(_3422_), .gnd(gnd), .vdd(vdd), .B(_3396_), .S(raddr1_4_bF_buf0_), );
  INVX1 INVX1_102 (.Y(_3423_), .A(regs_5__20_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1382 (.Y(_3424_), .A(_3423_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf78_), .C(raddr1_1_bF_buf11_bF_buf1_), );
  AOI21X1 AOI21X1_204 (.Y(_3425_), .A(regs_4__20_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf77_), .C(_3424_), );
  AND2X2 AND2X2_26 (.Y(_3426_), .A(regs_6__20_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf76_), );
  OAI21X1 OAI21X1_1383 (.Y(_3427_), .A(_2141_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf75_), .C(_2415__bF_buf6), );
  OAI21X1 OAI21X1_1384 (.Y(_3428_), .A(_3427_), .gnd(gnd), .vdd(vdd), .B(_3426_), .C(_2399__bF_buf5), );
  INVX1 INVX1_103 (.Y(_3429_), .A(regs_1__20_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1385 (.Y(_3430_), .A(_3429_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf74_), .C(raddr1_1_bF_buf10_bF_buf1_), );
  AOI21X1 AOI21X1_205 (.Y(_3431_), .A(regs_0__20_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf73_), .C(_3430_), );
  INVX1 INVX1_104 (.Y(_3432_), .A(regs_3__20_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_176 (.Y(_3433_), .A(raddr1_0_bF_buf72_), .gnd(gnd), .vdd(vdd), .B(_3432_), );
  NAND2X1 NAND2X1_549 (.Y(_3434_), .A(regs_2__20_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf71_), );
  NAND2X1 NAND2X1_550 (.Y(_3435_), .A(_2415__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_3434_), );
  OAI21X1 OAI21X1_1386 (.Y(_3436_), .A(_3435_), .gnd(gnd), .vdd(vdd), .B(_3433_), .C(raddr1_2_bF_buf3_), );
  OAI22X1 OAI22X1_34 (.Y(_3437_), .A(_3431_), .gnd(gnd), .vdd(vdd), .B(_3436_), .C(_3428_), .D(_3425_), );
  NAND2X1 NAND2X1_551 (.Y(_3438_), .A(regs_10__20_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf70_), );
  OAI21X1 OAI21X1_1387 (.Y(_3439_), .A(_1942_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf69_), .C(_3438_), );
  NAND2X1 NAND2X1_552 (.Y(_3440_), .A(regs_8__20_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf68_), );
  OAI21X1 OAI21X1_1388 (.Y(_3441_), .A(_2040_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf67_), .C(_3440_), );
  MUX2X1 MUX2X1_184 (.Y(_3442_), .A(_3441_), .gnd(gnd), .vdd(vdd), .B(_3439_), .S(raddr1_1_bF_buf9_bF_buf1_), );
  NAND2X1 NAND2X1_553 (.Y(_3443_), .A(regs_14__20_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf66_), );
  OAI21X1 OAI21X1_1389 (.Y(_3444_), .A(_1745_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf65_), .C(_3443_), );
  NAND2X1 NAND2X1_554 (.Y(_3445_), .A(regs_12__20_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf64_), );
  OAI21X1 OAI21X1_1390 (.Y(_3446_), .A(_1843_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf63_), .C(_3445_), );
  MUX2X1 MUX2X1_185 (.Y(_3447_), .A(_3446_), .gnd(gnd), .vdd(vdd), .B(_3444_), .S(raddr1_1_bF_buf8_), );
  MUX2X1 MUX2X1_186 (.Y(_3448_), .A(_3447_), .gnd(gnd), .vdd(vdd), .B(_3442_), .S(_2399__bF_buf4), );
  MUX2X1 MUX2X1_187 (.Y(_3449_), .A(_3448_), .gnd(gnd), .vdd(vdd), .B(_3437_), .S(_2398__bF_buf6), );
  OAI21X1 OAI21X1_1391 (.Y(_3450_), .A(_1645_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf62_), .C(raddr1_1_bF_buf7_), );
  AOI21X1 AOI21X1_206 (.Y(_3451_), .A(regs_16__20_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf61_), .C(_3450_), );
  NOR2X1 NOR2X1_177 (.Y(_3452_), .A(raddr1_0_bF_buf60_), .gnd(gnd), .vdd(vdd), .B(_1547_), );
  NAND2X1 NAND2X1_555 (.Y(_3453_), .A(regs_18__20_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf59_), );
  NAND2X1 NAND2X1_556 (.Y(_3454_), .A(_2415__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_3453_), );
  OAI21X1 OAI21X1_1392 (.Y(_3455_), .A(_3454_), .gnd(gnd), .vdd(vdd), .B(_3452_), .C(raddr1_2_bF_buf2_), );
  OAI21X1 OAI21X1_1393 (.Y(_3456_), .A(_1448_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf58_), .C(raddr1_1_bF_buf6_), );
  AOI21X1 AOI21X1_207 (.Y(_3457_), .A(regs_20__20_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf57_), .C(_3456_), );
  AND2X2 AND2X2_27 (.Y(_3458_), .A(regs_22__20_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf56_), );
  OAI21X1 OAI21X1_1394 (.Y(_3459_), .A(_1350_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf55_), .C(_2415__bF_buf3), );
  OAI21X1 OAI21X1_1395 (.Y(_3460_), .A(_3459_), .gnd(gnd), .vdd(vdd), .B(_3458_), .C(_2399__bF_buf3), );
  OAI22X1 OAI22X1_35 (.Y(_3461_), .A(_3451_), .gnd(gnd), .vdd(vdd), .B(_3455_), .C(_3460_), .D(_3457_), );
  INVX1 INVX1_105 (.Y(_3462_), .A(regs_29__20_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_557 (.Y(_3463_), .A(regs_28__20_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf54_), );
  OAI21X1 OAI21X1_1396 (.Y(_3464_), .A(_3462_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf53_), .C(_3463_), );
  MUX2X1 MUX2X1_188 (.Y(_3465_), .A(_3464_), .gnd(gnd), .vdd(vdd), .B(regs_30__20_), .S(raddr1_1_bF_buf5_), );
  NAND2X1 NAND2X1_558 (.Y(_3466_), .A(regs_26__20_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf52_), );
  OAI21X1 OAI21X1_1397 (.Y(_3467_), .A(_1183_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf51_), .C(_3466_), );
  INVX1 INVX1_106 (.Y(_3468_), .A(regs_25__20_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_559 (.Y(_3469_), .A(regs_24__20_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf50_), );
  OAI21X1 OAI21X1_1398 (.Y(_3470_), .A(_3468_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf49_), .C(_3469_), );
  MUX2X1 MUX2X1_189 (.Y(_3471_), .A(_3470_), .gnd(gnd), .vdd(vdd), .B(_3467_), .S(raddr1_1_bF_buf4_), );
  MUX2X1 MUX2X1_190 (.Y(_3472_), .A(_3471_), .gnd(gnd), .vdd(vdd), .B(_3465_), .S(raddr1_2_bF_buf1_), );
  MUX2X1 MUX2X1_191 (.Y(_3473_), .A(_3472_), .gnd(gnd), .vdd(vdd), .B(_3461_), .S(_2398__bF_buf5), );
  MUX2X1 MUX2X1_192 (.Y(_5511__20_), .A(_3449_), .gnd(gnd), .vdd(vdd), .B(_3473_), .S(raddr1_4_bF_buf4_), );
  INVX1 INVX1_107 (.Y(_3474_), .A(regs_5__21_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1399 (.Y(_3475_), .A(_3474_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf48_), .C(raddr1_1_bF_buf3_), );
  AOI21X1 AOI21X1_208 (.Y(_3476_), .A(regs_4__21_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf47_), .C(_3475_), );
  AND2X2 AND2X2_28 (.Y(_3477_), .A(regs_6__21_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf46_), );
  OAI21X1 OAI21X1_1400 (.Y(_3478_), .A(_2143_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf45_), .C(_2415__bF_buf2), );
  OAI21X1 OAI21X1_1401 (.Y(_3479_), .A(_3478_), .gnd(gnd), .vdd(vdd), .B(_3477_), .C(_2399__bF_buf2), );
  INVX1 INVX1_108 (.Y(_3480_), .A(regs_1__21_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1402 (.Y(_3481_), .A(_3480_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf44_), .C(raddr1_1_bF_buf2_), );
  AOI21X1 AOI21X1_209 (.Y(_3482_), .A(regs_0__21_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf43_), .C(_3481_), );
  INVX1 INVX1_109 (.Y(_3483_), .A(regs_3__21_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_178 (.Y(_3484_), .A(raddr1_0_bF_buf42_), .gnd(gnd), .vdd(vdd), .B(_3483_), );
  NAND2X1 NAND2X1_560 (.Y(_3485_), .A(regs_2__21_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf41_), );
  NAND2X1 NAND2X1_561 (.Y(_3486_), .A(_2415__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_3485_), );
  OAI21X1 OAI21X1_1403 (.Y(_3487_), .A(_3486_), .gnd(gnd), .vdd(vdd), .B(_3484_), .C(raddr1_2_bF_buf0_), );
  OAI22X1 OAI22X1_36 (.Y(_3488_), .A(_3482_), .gnd(gnd), .vdd(vdd), .B(_3487_), .C(_3479_), .D(_3476_), );
  NAND2X1 NAND2X1_562 (.Y(_3489_), .A(regs_10__21_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf40_), );
  OAI21X1 OAI21X1_1404 (.Y(_3490_), .A(_1944_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf39_), .C(_3489_), );
  NAND2X1 NAND2X1_563 (.Y(_3491_), .A(regs_8__21_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf38_), );
  OAI21X1 OAI21X1_1405 (.Y(_3492_), .A(_2042_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf37_), .C(_3491_), );
  MUX2X1 MUX2X1_193 (.Y(_3493_), .A(_3492_), .gnd(gnd), .vdd(vdd), .B(_3490_), .S(raddr1_1_bF_buf1_), );
  NAND2X1 NAND2X1_564 (.Y(_3494_), .A(regs_14__21_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf36_), );
  OAI21X1 OAI21X1_1406 (.Y(_3495_), .A(_1747_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf35_), .C(_3494_), );
  NAND2X1 NAND2X1_565 (.Y(_3496_), .A(regs_12__21_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf34_), );
  OAI21X1 OAI21X1_1407 (.Y(_3497_), .A(_1845_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf33_), .C(_3496_), );
  MUX2X1 MUX2X1_194 (.Y(_3498_), .A(_3497_), .gnd(gnd), .vdd(vdd), .B(_3495_), .S(raddr1_1_bF_buf0_), );
  MUX2X1 MUX2X1_195 (.Y(_3499_), .A(_3498_), .gnd(gnd), .vdd(vdd), .B(_3493_), .S(_2399__bF_buf1), );
  MUX2X1 MUX2X1_196 (.Y(_3500_), .A(_3499_), .gnd(gnd), .vdd(vdd), .B(_3488_), .S(_2398__bF_buf4), );
  OAI21X1 OAI21X1_1408 (.Y(_3501_), .A(_1647_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf32_), .C(raddr1_1_bF_buf14_bF_buf0_), );
  AOI21X1 AOI21X1_210 (.Y(_3502_), .A(regs_16__21_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf31_), .C(_3501_), );
  NOR2X1 NOR2X1_179 (.Y(_3503_), .A(raddr1_0_bF_buf30_), .gnd(gnd), .vdd(vdd), .B(_1549_), );
  NAND2X1 NAND2X1_566 (.Y(_3504_), .A(regs_18__21_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf29_), );
  NAND2X1 NAND2X1_567 (.Y(_3505_), .A(_2415__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_3504_), );
  OAI21X1 OAI21X1_1409 (.Y(_3506_), .A(_3505_), .gnd(gnd), .vdd(vdd), .B(_3503_), .C(raddr1_2_bF_buf10_), );
  OAI21X1 OAI21X1_1410 (.Y(_3507_), .A(_1450_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf28_), .C(raddr1_1_bF_buf13_bF_buf0_), );
  AOI21X1 AOI21X1_211 (.Y(_3508_), .A(regs_20__21_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf27_), .C(_3507_), );
  AND2X2 AND2X2_29 (.Y(_3509_), .A(regs_22__21_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf26_), );
  OAI21X1 OAI21X1_1411 (.Y(_3510_), .A(_1352_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf25_), .C(_2415__bF_buf8), );
  OAI21X1 OAI21X1_1412 (.Y(_3511_), .A(_3510_), .gnd(gnd), .vdd(vdd), .B(_3509_), .C(_2399__bF_buf0), );
  OAI22X1 OAI22X1_37 (.Y(_3512_), .A(_3502_), .gnd(gnd), .vdd(vdd), .B(_3506_), .C(_3511_), .D(_3508_), );
  INVX1 INVX1_110 (.Y(_3513_), .A(regs_29__21_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_568 (.Y(_3514_), .A(regs_28__21_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf24_), );
  OAI21X1 OAI21X1_1413 (.Y(_3515_), .A(_3513_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf23_), .C(_3514_), );
  MUX2X1 MUX2X1_197 (.Y(_3516_), .A(_3515_), .gnd(gnd), .vdd(vdd), .B(regs_30__21_), .S(raddr1_1_bF_buf12_bF_buf0_), );
  NAND2X1 NAND2X1_569 (.Y(_3517_), .A(regs_26__21_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf22_), );
  OAI21X1 OAI21X1_1414 (.Y(_3518_), .A(_1185_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf21_), .C(_3517_), );
  INVX1 INVX1_111 (.Y(_3519_), .A(regs_25__21_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_570 (.Y(_3520_), .A(regs_24__21_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf20_), );
  OAI21X1 OAI21X1_1415 (.Y(_3521_), .A(_3519_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf19_), .C(_3520_), );
  MUX2X1 MUX2X1_198 (.Y(_3522_), .A(_3521_), .gnd(gnd), .vdd(vdd), .B(_3518_), .S(raddr1_1_bF_buf11_bF_buf0_), );
  MUX2X1 MUX2X1_199 (.Y(_3523_), .A(_3522_), .gnd(gnd), .vdd(vdd), .B(_3516_), .S(raddr1_2_bF_buf9_), );
  MUX2X1 MUX2X1_200 (.Y(_3524_), .A(_3523_), .gnd(gnd), .vdd(vdd), .B(_3512_), .S(_2398__bF_buf3), );
  MUX2X1 MUX2X1_201 (.Y(_5511__21_), .A(_3500_), .gnd(gnd), .vdd(vdd), .B(_3524_), .S(raddr1_4_bF_buf3_), );
  OAI21X1 OAI21X1_1416 (.Y(_3525_), .A(_1452_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf18_), .C(raddr1_1_bF_buf10_bF_buf0_), );
  AOI21X1 AOI21X1_212 (.Y(_3526_), .A(regs_20__22_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf17_), .C(_3525_), );
  AND2X2 AND2X2_30 (.Y(_3527_), .A(regs_22__22_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf16_), );
  OAI21X1 OAI21X1_1417 (.Y(_3528_), .A(_1354_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf15_), .C(_2415__bF_buf7), );
  OAI21X1 OAI21X1_1418 (.Y(_3529_), .A(_3528_), .gnd(gnd), .vdd(vdd), .B(_3527_), .C(_2399__bF_buf8), );
  OAI21X1 OAI21X1_1419 (.Y(_3530_), .A(_1649_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf14_), .C(raddr1_1_bF_buf9_bF_buf0_), );
  AOI21X1 AOI21X1_213 (.Y(_3531_), .A(regs_16__22_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf13_), .C(_3530_), );
  NOR2X1 NOR2X1_180 (.Y(_3532_), .A(raddr1_0_bF_buf12_), .gnd(gnd), .vdd(vdd), .B(_1551_), );
  NAND2X1 NAND2X1_571 (.Y(_3533_), .A(regs_18__22_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf11_), );
  NAND2X1 NAND2X1_572 (.Y(_3534_), .A(_2415__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_3533_), );
  OAI21X1 OAI21X1_1420 (.Y(_3535_), .A(_3534_), .gnd(gnd), .vdd(vdd), .B(_3532_), .C(raddr1_2_bF_buf8_), );
  OAI22X1 OAI22X1_38 (.Y(_3536_), .A(_3531_), .gnd(gnd), .vdd(vdd), .B(_3535_), .C(_3529_), .D(_3526_), );
  INVX1 INVX1_112 (.Y(_3537_), .A(regs_29__22_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_573 (.Y(_3538_), .A(regs_28__22_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf10_), );
  OAI21X1 OAI21X1_1421 (.Y(_3539_), .A(_3537_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf9_), .C(_3538_), );
  MUX2X1 MUX2X1_202 (.Y(_3540_), .A(_3539_), .gnd(gnd), .vdd(vdd), .B(regs_30__22_), .S(raddr1_1_bF_buf8_), );
  NAND2X1 NAND2X1_574 (.Y(_3541_), .A(regs_26__22_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf8_), );
  OAI21X1 OAI21X1_1422 (.Y(_3542_), .A(_1187_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf7_), .C(_3541_), );
  INVX1 INVX1_113 (.Y(_3543_), .A(regs_25__22_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_575 (.Y(_3544_), .A(regs_24__22_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf6_), );
  OAI21X1 OAI21X1_1423 (.Y(_3545_), .A(_3543_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf5_), .C(_3544_), );
  MUX2X1 MUX2X1_203 (.Y(_3546_), .A(_3545_), .gnd(gnd), .vdd(vdd), .B(_3542_), .S(raddr1_1_bF_buf7_), );
  MUX2X1 MUX2X1_204 (.Y(_3547_), .A(_3546_), .gnd(gnd), .vdd(vdd), .B(_3540_), .S(raddr1_2_bF_buf7_), );
  MUX2X1 MUX2X1_205 (.Y(_3548_), .A(_3547_), .gnd(gnd), .vdd(vdd), .B(_3536_), .S(_2398__bF_buf2), );
  NAND2X1 NAND2X1_576 (.Y(_3549_), .A(regs_6__22_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf4_), );
  OAI21X1 OAI21X1_1424 (.Y(_3550_), .A(_2145_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf3_), .C(_3549_), );
  INVX1 INVX1_114 (.Y(_3551_), .A(regs_5__22_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_577 (.Y(_3552_), .A(regs_4__22_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf2_), );
  OAI21X1 OAI21X1_1425 (.Y(_3553_), .A(_3551_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf1_), .C(_3552_), );
  MUX2X1 MUX2X1_206 (.Y(_3554_), .A(_3553_), .gnd(gnd), .vdd(vdd), .B(_3550_), .S(raddr1_1_bF_buf6_), );
  INVX1 INVX1_115 (.Y(_3555_), .A(regs_3__22_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_578 (.Y(_3556_), .A(regs_2__22_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf0_), );
  OAI21X1 OAI21X1_1426 (.Y(_3557_), .A(_3555_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf96_), .C(_3556_), );
  INVX1 INVX1_116 (.Y(_3558_), .A(regs_1__22_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_579 (.Y(_3559_), .A(regs_0__22_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf95_), );
  OAI21X1 OAI21X1_1427 (.Y(_3560_), .A(_3558_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf94_), .C(_3559_), );
  MUX2X1 MUX2X1_207 (.Y(_3561_), .A(_3560_), .gnd(gnd), .vdd(vdd), .B(_3557_), .S(raddr1_1_bF_buf5_), );
  MUX2X1 MUX2X1_208 (.Y(_3562_), .A(_3561_), .gnd(gnd), .vdd(vdd), .B(_3554_), .S(raddr1_2_bF_buf6_), );
  NAND2X1 NAND2X1_580 (.Y(_3563_), .A(regs_14__22_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf93_), );
  OAI21X1 OAI21X1_1428 (.Y(_3564_), .A(_1749_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf92_), .C(_3563_), );
  NAND2X1 NAND2X1_581 (.Y(_3565_), .A(regs_12__22_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf91_), );
  OAI21X1 OAI21X1_1429 (.Y(_3566_), .A(_1847_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf90_), .C(_3565_), );
  MUX2X1 MUX2X1_209 (.Y(_3567_), .A(_3566_), .gnd(gnd), .vdd(vdd), .B(_3564_), .S(raddr1_1_bF_buf4_), );
  NAND2X1 NAND2X1_582 (.Y(_3568_), .A(regs_10__22_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf89_), );
  OAI21X1 OAI21X1_1430 (.Y(_3569_), .A(_1946_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf88_), .C(_3568_), );
  NAND2X1 NAND2X1_583 (.Y(_3570_), .A(regs_8__22_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf87_), );
  OAI21X1 OAI21X1_1431 (.Y(_3571_), .A(_2044_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf86_), .C(_3570_), );
  MUX2X1 MUX2X1_210 (.Y(_3572_), .A(_3571_), .gnd(gnd), .vdd(vdd), .B(_3569_), .S(raddr1_1_bF_buf3_), );
  MUX2X1 MUX2X1_211 (.Y(_3573_), .A(_3572_), .gnd(gnd), .vdd(vdd), .B(_3567_), .S(raddr1_2_bF_buf5_), );
  MUX2X1 MUX2X1_212 (.Y(_3574_), .A(_3573_), .gnd(gnd), .vdd(vdd), .B(_3562_), .S(_2398__bF_buf1), );
  MUX2X1 MUX2X1_213 (.Y(_5511__22_), .A(_3574_), .gnd(gnd), .vdd(vdd), .B(_3548_), .S(raddr1_4_bF_buf2_), );
  OAI21X1 OAI21X1_1432 (.Y(_3575_), .A(_1454_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf85_), .C(raddr1_1_bF_buf2_), );
  AOI21X1 AOI21X1_214 (.Y(_3576_), .A(regs_20__23_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf84_), .C(_3575_), );
  AND2X2 AND2X2_31 (.Y(_3577_), .A(regs_22__23_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf83_), );
  OAI21X1 OAI21X1_1433 (.Y(_3578_), .A(_1356_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf82_), .C(_2415__bF_buf5), );
  OAI21X1 OAI21X1_1434 (.Y(_3579_), .A(_3578_), .gnd(gnd), .vdd(vdd), .B(_3577_), .C(_2399__bF_buf7), );
  OAI21X1 OAI21X1_1435 (.Y(_3580_), .A(_1651_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf81_), .C(raddr1_1_bF_buf1_), );
  AOI21X1 AOI21X1_215 (.Y(_3581_), .A(regs_16__23_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf80_), .C(_3580_), );
  NOR2X1 NOR2X1_181 (.Y(_3582_), .A(raddr1_0_bF_buf79_), .gnd(gnd), .vdd(vdd), .B(_1553_), );
  NAND2X1 NAND2X1_584 (.Y(_3583_), .A(regs_18__23_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf78_), );
  NAND2X1 NAND2X1_585 (.Y(_3584_), .A(_2415__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_3583_), );
  OAI21X1 OAI21X1_1436 (.Y(_3585_), .A(_3584_), .gnd(gnd), .vdd(vdd), .B(_3582_), .C(raddr1_2_bF_buf4_), );
  OAI22X1 OAI22X1_39 (.Y(_3586_), .A(_3581_), .gnd(gnd), .vdd(vdd), .B(_3585_), .C(_3579_), .D(_3576_), );
  INVX1 INVX1_117 (.Y(_3587_), .A(regs_29__23_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_586 (.Y(_3588_), .A(regs_28__23_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf77_), );
  OAI21X1 OAI21X1_1437 (.Y(_3589_), .A(_3587_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf76_), .C(_3588_), );
  MUX2X1 MUX2X1_214 (.Y(_3590_), .A(_3589_), .gnd(gnd), .vdd(vdd), .B(regs_30__23_), .S(raddr1_1_bF_buf0_), );
  NAND2X1 NAND2X1_587 (.Y(_3591_), .A(regs_26__23_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf75_), );
  OAI21X1 OAI21X1_1438 (.Y(_3592_), .A(_1189_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf74_), .C(_3591_), );
  INVX1 INVX1_118 (.Y(_3593_), .A(regs_25__23_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_588 (.Y(_3594_), .A(regs_24__23_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf73_), );
  OAI21X1 OAI21X1_1439 (.Y(_3595_), .A(_3593_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf72_), .C(_3594_), );
  MUX2X1 MUX2X1_215 (.Y(_3596_), .A(_3595_), .gnd(gnd), .vdd(vdd), .B(_3592_), .S(raddr1_1_bF_buf14_bF_buf3_), );
  MUX2X1 MUX2X1_216 (.Y(_3597_), .A(_3596_), .gnd(gnd), .vdd(vdd), .B(_3590_), .S(raddr1_2_bF_buf3_), );
  MUX2X1 MUX2X1_217 (.Y(_3598_), .A(_3597_), .gnd(gnd), .vdd(vdd), .B(_3586_), .S(_2398__bF_buf0), );
  NAND2X1 NAND2X1_589 (.Y(_3599_), .A(regs_6__23_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf71_), );
  OAI21X1 OAI21X1_1440 (.Y(_3600_), .A(_2147_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf70_), .C(_3599_), );
  INVX1 INVX1_119 (.Y(_3601_), .A(regs_5__23_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_590 (.Y(_3602_), .A(regs_4__23_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf69_), );
  OAI21X1 OAI21X1_1441 (.Y(_3603_), .A(_3601_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf68_), .C(_3602_), );
  MUX2X1 MUX2X1_218 (.Y(_3604_), .A(_3603_), .gnd(gnd), .vdd(vdd), .B(_3600_), .S(raddr1_1_bF_buf13_bF_buf3_), );
  INVX1 INVX1_120 (.Y(_3605_), .A(regs_3__23_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_591 (.Y(_3606_), .A(regs_2__23_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf67_), );
  OAI21X1 OAI21X1_1442 (.Y(_3607_), .A(_3605_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf66_), .C(_3606_), );
  INVX1 INVX1_121 (.Y(_3608_), .A(regs_1__23_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_592 (.Y(_3609_), .A(regs_0__23_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf65_), );
  OAI21X1 OAI21X1_1443 (.Y(_3610_), .A(_3608_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf64_), .C(_3609_), );
  MUX2X1 MUX2X1_219 (.Y(_3611_), .A(_3610_), .gnd(gnd), .vdd(vdd), .B(_3607_), .S(raddr1_1_bF_buf12_bF_buf3_), );
  MUX2X1 MUX2X1_220 (.Y(_3612_), .A(_3611_), .gnd(gnd), .vdd(vdd), .B(_3604_), .S(raddr1_2_bF_buf2_), );
  NAND2X1 NAND2X1_593 (.Y(_3613_), .A(regs_14__23_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf63_), );
  OAI21X1 OAI21X1_1444 (.Y(_3614_), .A(_1751_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf62_), .C(_3613_), );
  NAND2X1 NAND2X1_594 (.Y(_3615_), .A(regs_12__23_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf61_), );
  OAI21X1 OAI21X1_1445 (.Y(_3616_), .A(_1849_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf60_), .C(_3615_), );
  MUX2X1 MUX2X1_221 (.Y(_3617_), .A(_3616_), .gnd(gnd), .vdd(vdd), .B(_3614_), .S(raddr1_1_bF_buf11_bF_buf3_), );
  NAND2X1 NAND2X1_595 (.Y(_3618_), .A(regs_10__23_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf59_), );
  OAI21X1 OAI21X1_1446 (.Y(_3619_), .A(_1948_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf58_), .C(_3618_), );
  NAND2X1 NAND2X1_596 (.Y(_3620_), .A(regs_8__23_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf57_), );
  OAI21X1 OAI21X1_1447 (.Y(_3621_), .A(_2046_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf56_), .C(_3620_), );
  MUX2X1 MUX2X1_222 (.Y(_3622_), .A(_3621_), .gnd(gnd), .vdd(vdd), .B(_3619_), .S(raddr1_1_bF_buf10_bF_buf3_), );
  MUX2X1 MUX2X1_223 (.Y(_3623_), .A(_3622_), .gnd(gnd), .vdd(vdd), .B(_3617_), .S(raddr1_2_bF_buf1_), );
  MUX2X1 MUX2X1_224 (.Y(_3624_), .A(_3623_), .gnd(gnd), .vdd(vdd), .B(_3612_), .S(_2398__bF_buf7), );
  MUX2X1 MUX2X1_225 (.Y(_5511__23_), .A(_3624_), .gnd(gnd), .vdd(vdd), .B(_3598_), .S(raddr1_4_bF_buf1_), );
  OAI21X1 OAI21X1_1448 (.Y(_3625_), .A(_1456_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf55_), .C(raddr1_1_bF_buf9_bF_buf3_), );
  AOI21X1 AOI21X1_216 (.Y(_3626_), .A(regs_20__24_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf54_), .C(_3625_), );
  AND2X2 AND2X2_32 (.Y(_3627_), .A(regs_22__24_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf53_), );
  OAI21X1 OAI21X1_1449 (.Y(_3628_), .A(_1358_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf52_), .C(_2415__bF_buf3), );
  OAI21X1 OAI21X1_1450 (.Y(_3629_), .A(_3628_), .gnd(gnd), .vdd(vdd), .B(_3627_), .C(_2399__bF_buf6), );
  OAI21X1 OAI21X1_1451 (.Y(_3630_), .A(_1653_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf51_), .C(raddr1_1_bF_buf8_), );
  AOI21X1 AOI21X1_217 (.Y(_3631_), .A(regs_16__24_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf50_), .C(_3630_), );
  NOR2X1 NOR2X1_182 (.Y(_3632_), .A(raddr1_0_bF_buf49_), .gnd(gnd), .vdd(vdd), .B(_1555_), );
  NAND2X1 NAND2X1_597 (.Y(_3633_), .A(regs_18__24_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf48_), );
  NAND2X1 NAND2X1_598 (.Y(_3634_), .A(_2415__bF_buf2), .gnd(gnd), .vdd(vdd), .B(_3633_), );
  OAI21X1 OAI21X1_1452 (.Y(_3635_), .A(_3634_), .gnd(gnd), .vdd(vdd), .B(_3632_), .C(raddr1_2_bF_buf0_), );
  OAI22X1 OAI22X1_40 (.Y(_3636_), .A(_3631_), .gnd(gnd), .vdd(vdd), .B(_3635_), .C(_3629_), .D(_3626_), );
  INVX1 INVX1_122 (.Y(_3637_), .A(regs_29__24_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_599 (.Y(_3638_), .A(regs_28__24_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf47_), );
  OAI21X1 OAI21X1_1453 (.Y(_3639_), .A(_3637_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf46_), .C(_3638_), );
  MUX2X1 MUX2X1_226 (.Y(_3640_), .A(_3639_), .gnd(gnd), .vdd(vdd), .B(regs_30__24_), .S(raddr1_1_bF_buf7_), );
  NAND2X1 NAND2X1_600 (.Y(_3641_), .A(regs_26__24_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf45_), );
  OAI21X1 OAI21X1_1454 (.Y(_3642_), .A(_1191_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf44_), .C(_3641_), );
  INVX1 INVX1_123 (.Y(_3643_), .A(regs_25__24_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_601 (.Y(_3644_), .A(regs_24__24_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf43_), );
  OAI21X1 OAI21X1_1455 (.Y(_3645_), .A(_3643_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf42_), .C(_3644_), );
  MUX2X1 MUX2X1_227 (.Y(_3646_), .A(_3645_), .gnd(gnd), .vdd(vdd), .B(_3642_), .S(raddr1_1_bF_buf6_), );
  MUX2X1 MUX2X1_228 (.Y(_3647_), .A(_3646_), .gnd(gnd), .vdd(vdd), .B(_3640_), .S(raddr1_2_bF_buf10_), );
  MUX2X1 MUX2X1_229 (.Y(_3648_), .A(_3647_), .gnd(gnd), .vdd(vdd), .B(_3636_), .S(_2398__bF_buf6), );
  NAND2X1 NAND2X1_602 (.Y(_3649_), .A(regs_6__24_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf41_), );
  OAI21X1 OAI21X1_1456 (.Y(_3650_), .A(_2149_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf40_), .C(_3649_), );
  INVX1 INVX1_124 (.Y(_3651_), .A(regs_5__24_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_603 (.Y(_3652_), .A(regs_4__24_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf39_), );
  OAI21X1 OAI21X1_1457 (.Y(_3653_), .A(_3651_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf38_), .C(_3652_), );
  MUX2X1 MUX2X1_230 (.Y(_3654_), .A(_3653_), .gnd(gnd), .vdd(vdd), .B(_3650_), .S(raddr1_1_bF_buf5_), );
  INVX1 INVX1_125 (.Y(_3655_), .A(regs_3__24_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_604 (.Y(_3656_), .A(regs_2__24_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf37_), );
  OAI21X1 OAI21X1_1458 (.Y(_3657_), .A(_3655_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf36_), .C(_3656_), );
  INVX1 INVX1_126 (.Y(_3658_), .A(regs_1__24_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_605 (.Y(_3659_), .A(regs_0__24_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf35_), );
  OAI21X1 OAI21X1_1459 (.Y(_3660_), .A(_3658_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf34_), .C(_3659_), );
  MUX2X1 MUX2X1_231 (.Y(_3661_), .A(_3660_), .gnd(gnd), .vdd(vdd), .B(_3657_), .S(raddr1_1_bF_buf4_), );
  MUX2X1 MUX2X1_232 (.Y(_3662_), .A(_3661_), .gnd(gnd), .vdd(vdd), .B(_3654_), .S(raddr1_2_bF_buf9_), );
  NAND2X1 NAND2X1_606 (.Y(_3663_), .A(regs_10__24_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf33_), );
  OAI21X1 OAI21X1_1460 (.Y(_3664_), .A(_1950_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf32_), .C(_3663_), );
  NAND2X1 NAND2X1_607 (.Y(_3665_), .A(regs_8__24_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf31_), );
  OAI21X1 OAI21X1_1461 (.Y(_3666_), .A(_2048_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf30_), .C(_3665_), );
  MUX2X1 MUX2X1_233 (.Y(_3667_), .A(_3666_), .gnd(gnd), .vdd(vdd), .B(_3664_), .S(raddr1_1_bF_buf3_), );
  NAND2X1 NAND2X1_608 (.Y(_3668_), .A(regs_14__24_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf29_), );
  OAI21X1 OAI21X1_1462 (.Y(_3669_), .A(_1753_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf28_), .C(_3668_), );
  NAND2X1 NAND2X1_609 (.Y(_3670_), .A(regs_12__24_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf27_), );
  OAI21X1 OAI21X1_1463 (.Y(_3671_), .A(_1851_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf26_), .C(_3670_), );
  MUX2X1 MUX2X1_234 (.Y(_3672_), .A(_3671_), .gnd(gnd), .vdd(vdd), .B(_3669_), .S(raddr1_1_bF_buf2_), );
  MUX2X1 MUX2X1_235 (.Y(_3673_), .A(_3672_), .gnd(gnd), .vdd(vdd), .B(_3667_), .S(_2399__bF_buf5), );
  MUX2X1 MUX2X1_236 (.Y(_3674_), .A(_3673_), .gnd(gnd), .vdd(vdd), .B(_3662_), .S(_2398__bF_buf5), );
  MUX2X1 MUX2X1_237 (.Y(_5511__24_), .A(_3674_), .gnd(gnd), .vdd(vdd), .B(_3648_), .S(raddr1_4_bF_buf0_), );
  INVX1 INVX1_127 (.Y(_3675_), .A(regs_5__25_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1464 (.Y(_3676_), .A(_3675_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf25_), .C(raddr1_1_bF_buf1_), );
  AOI21X1 AOI21X1_218 (.Y(_3677_), .A(regs_4__25_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf24_), .C(_3676_), );
  AND2X2 AND2X2_33 (.Y(_3678_), .A(regs_6__25_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf23_), );
  OAI21X1 OAI21X1_1465 (.Y(_3679_), .A(_2151_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf22_), .C(_2415__bF_buf1), );
  OAI21X1 OAI21X1_1466 (.Y(_3680_), .A(_3679_), .gnd(gnd), .vdd(vdd), .B(_3678_), .C(_2399__bF_buf4), );
  INVX1 INVX1_128 (.Y(_3681_), .A(regs_1__25_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1467 (.Y(_3682_), .A(_3681_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf21_), .C(raddr1_1_bF_buf0_), );
  AOI21X1 AOI21X1_219 (.Y(_3683_), .A(regs_0__25_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf20_), .C(_3682_), );
  INVX1 INVX1_129 (.Y(_3684_), .A(regs_3__25_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_183 (.Y(_3685_), .A(raddr1_0_bF_buf19_), .gnd(gnd), .vdd(vdd), .B(_3684_), );
  NAND2X1 NAND2X1_610 (.Y(_3686_), .A(regs_2__25_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf18_), );
  NAND2X1 NAND2X1_611 (.Y(_3687_), .A(_2415__bF_buf0), .gnd(gnd), .vdd(vdd), .B(_3686_), );
  OAI21X1 OAI21X1_1468 (.Y(_3688_), .A(_3687_), .gnd(gnd), .vdd(vdd), .B(_3685_), .C(raddr1_2_bF_buf8_), );
  OAI22X1 OAI22X1_41 (.Y(_3689_), .A(_3683_), .gnd(gnd), .vdd(vdd), .B(_3688_), .C(_3680_), .D(_3677_), );
  NAND2X1 NAND2X1_612 (.Y(_3690_), .A(regs_10__25_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf17_), );
  OAI21X1 OAI21X1_1469 (.Y(_3691_), .A(_1952_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf16_), .C(_3690_), );
  NAND2X1 NAND2X1_613 (.Y(_3692_), .A(regs_8__25_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf15_), );
  OAI21X1 OAI21X1_1470 (.Y(_3693_), .A(_2050_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf14_), .C(_3692_), );
  MUX2X1 MUX2X1_238 (.Y(_3694_), .A(_3693_), .gnd(gnd), .vdd(vdd), .B(_3691_), .S(raddr1_1_bF_buf14_bF_buf2_), );
  NAND2X1 NAND2X1_614 (.Y(_3695_), .A(regs_14__25_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf13_), );
  OAI21X1 OAI21X1_1471 (.Y(_3696_), .A(_1755_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf12_), .C(_3695_), );
  NAND2X1 NAND2X1_615 (.Y(_3697_), .A(regs_12__25_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf11_), );
  OAI21X1 OAI21X1_1472 (.Y(_3698_), .A(_1853_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf10_), .C(_3697_), );
  MUX2X1 MUX2X1_239 (.Y(_3699_), .A(_3698_), .gnd(gnd), .vdd(vdd), .B(_3696_), .S(raddr1_1_bF_buf13_bF_buf2_), );
  MUX2X1 MUX2X1_240 (.Y(_3700_), .A(_3699_), .gnd(gnd), .vdd(vdd), .B(_3694_), .S(_2399__bF_buf3), );
  MUX2X1 MUX2X1_241 (.Y(_3701_), .A(_3700_), .gnd(gnd), .vdd(vdd), .B(_3689_), .S(_2398__bF_buf4), );
  OAI21X1 OAI21X1_1473 (.Y(_3702_), .A(_1655_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf9_), .C(raddr1_1_bF_buf12_bF_buf2_), );
  AOI21X1 AOI21X1_220 (.Y(_3703_), .A(regs_16__25_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf8_), .C(_3702_), );
  NOR2X1 NOR2X1_184 (.Y(_3704_), .A(raddr1_0_bF_buf7_), .gnd(gnd), .vdd(vdd), .B(_1557_), );
  NAND2X1 NAND2X1_616 (.Y(_3705_), .A(regs_18__25_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf6_), );
  NAND2X1 NAND2X1_617 (.Y(_3706_), .A(_2415__bF_buf8), .gnd(gnd), .vdd(vdd), .B(_3705_), );
  OAI21X1 OAI21X1_1474 (.Y(_3707_), .A(_3706_), .gnd(gnd), .vdd(vdd), .B(_3704_), .C(raddr1_2_bF_buf7_), );
  OAI21X1 OAI21X1_1475 (.Y(_3708_), .A(_1458_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf5_), .C(raddr1_1_bF_buf11_bF_buf2_), );
  AOI21X1 AOI21X1_221 (.Y(_3709_), .A(regs_20__25_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf4_), .C(_3708_), );
  AND2X2 AND2X2_34 (.Y(_3710_), .A(regs_22__25_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf3_), );
  OAI21X1 OAI21X1_1476 (.Y(_3711_), .A(_1360_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf2_), .C(_2415__bF_buf7), );
  OAI21X1 OAI21X1_1477 (.Y(_3712_), .A(_3711_), .gnd(gnd), .vdd(vdd), .B(_3710_), .C(_2399__bF_buf2), );
  OAI22X1 OAI22X1_42 (.Y(_3713_), .A(_3703_), .gnd(gnd), .vdd(vdd), .B(_3707_), .C(_3712_), .D(_3709_), );
  INVX1 INVX1_130 (.Y(_3714_), .A(regs_29__25_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_618 (.Y(_3715_), .A(regs_28__25_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf1_), );
  OAI21X1 OAI21X1_1478 (.Y(_3716_), .A(_3714_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf0_), .C(_3715_), );
  MUX2X1 MUX2X1_242 (.Y(_3717_), .A(_3716_), .gnd(gnd), .vdd(vdd), .B(regs_30__25_), .S(raddr1_1_bF_buf10_bF_buf2_), );
  NAND2X1 NAND2X1_619 (.Y(_3718_), .A(regs_26__25_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf96_), );
  OAI21X1 OAI21X1_1479 (.Y(_3719_), .A(_1193_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf95_), .C(_3718_), );
  INVX1 INVX1_131 (.Y(_3720_), .A(regs_25__25_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_620 (.Y(_3721_), .A(regs_24__25_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf94_), );
  OAI21X1 OAI21X1_1480 (.Y(_3722_), .A(_3720_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf93_), .C(_3721_), );
  MUX2X1 MUX2X1_243 (.Y(_3723_), .A(_3722_), .gnd(gnd), .vdd(vdd), .B(_3719_), .S(raddr1_1_bF_buf9_bF_buf2_), );
  MUX2X1 MUX2X1_244 (.Y(_3724_), .A(_3723_), .gnd(gnd), .vdd(vdd), .B(_3717_), .S(raddr1_2_bF_buf6_), );
  MUX2X1 MUX2X1_245 (.Y(_3725_), .A(_3724_), .gnd(gnd), .vdd(vdd), .B(_3713_), .S(_2398__bF_buf3), );
  MUX2X1 MUX2X1_246 (.Y(_5511__25_), .A(_3701_), .gnd(gnd), .vdd(vdd), .B(_3725_), .S(raddr1_4_bF_buf4_), );
  INVX1 INVX1_132 (.Y(_3726_), .A(regs_5__26_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1481 (.Y(_3727_), .A(_3726_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf92_), .C(raddr1_1_bF_buf8_), );
  AOI21X1 AOI21X1_222 (.Y(_3728_), .A(regs_4__26_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf91_), .C(_3727_), );
  AND2X2 AND2X2_35 (.Y(_3729_), .A(regs_6__26_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf90_), );
  OAI21X1 OAI21X1_1482 (.Y(_3730_), .A(_2153_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf89_), .C(_2415__bF_buf6), );
  OAI21X1 OAI21X1_1483 (.Y(_3731_), .A(_3730_), .gnd(gnd), .vdd(vdd), .B(_3729_), .C(_2399__bF_buf1), );
  INVX1 INVX1_133 (.Y(_3732_), .A(regs_1__26_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1484 (.Y(_3733_), .A(_3732_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf88_), .C(raddr1_1_bF_buf7_), );
  AOI21X1 AOI21X1_223 (.Y(_3734_), .A(regs_0__26_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf87_), .C(_3733_), );
  INVX1 INVX1_134 (.Y(_3735_), .A(regs_3__26_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_185 (.Y(_3736_), .A(raddr1_0_bF_buf86_), .gnd(gnd), .vdd(vdd), .B(_3735_), );
  NAND2X1 NAND2X1_621 (.Y(_3737_), .A(regs_2__26_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf85_), );
  NAND2X1 NAND2X1_622 (.Y(_3738_), .A(_2415__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_3737_), );
  OAI21X1 OAI21X1_1485 (.Y(_3739_), .A(_3738_), .gnd(gnd), .vdd(vdd), .B(_3736_), .C(raddr1_2_bF_buf5_), );
  OAI22X1 OAI22X1_43 (.Y(_3740_), .A(_3734_), .gnd(gnd), .vdd(vdd), .B(_3739_), .C(_3731_), .D(_3728_), );
  NAND2X1 NAND2X1_623 (.Y(_3741_), .A(regs_10__26_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf84_), );
  OAI21X1 OAI21X1_1486 (.Y(_3742_), .A(_1954_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf83_), .C(_3741_), );
  NAND2X1 NAND2X1_624 (.Y(_3743_), .A(regs_8__26_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf82_), );
  OAI21X1 OAI21X1_1487 (.Y(_3744_), .A(_2052_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf81_), .C(_3743_), );
  MUX2X1 MUX2X1_247 (.Y(_3745_), .A(_3744_), .gnd(gnd), .vdd(vdd), .B(_3742_), .S(raddr1_1_bF_buf6_), );
  NAND2X1 NAND2X1_625 (.Y(_3746_), .A(regs_14__26_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf80_), );
  OAI21X1 OAI21X1_1488 (.Y(_3747_), .A(_1757_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf79_), .C(_3746_), );
  NAND2X1 NAND2X1_626 (.Y(_3748_), .A(regs_12__26_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf78_), );
  OAI21X1 OAI21X1_1489 (.Y(_3749_), .A(_1855_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf77_), .C(_3748_), );
  MUX2X1 MUX2X1_248 (.Y(_3750_), .A(_3749_), .gnd(gnd), .vdd(vdd), .B(_3747_), .S(raddr1_1_bF_buf5_), );
  MUX2X1 MUX2X1_249 (.Y(_3751_), .A(_3750_), .gnd(gnd), .vdd(vdd), .B(_3745_), .S(_2399__bF_buf0), );
  MUX2X1 MUX2X1_250 (.Y(_3752_), .A(_3751_), .gnd(gnd), .vdd(vdd), .B(_3740_), .S(_2398__bF_buf2), );
  OAI21X1 OAI21X1_1490 (.Y(_3753_), .A(_1657_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf76_), .C(raddr1_1_bF_buf4_), );
  AOI21X1 AOI21X1_224 (.Y(_3754_), .A(regs_16__26_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf75_), .C(_3753_), );
  NOR2X1 NOR2X1_186 (.Y(_3755_), .A(raddr1_0_bF_buf74_), .gnd(gnd), .vdd(vdd), .B(_1559_), );
  NAND2X1 NAND2X1_627 (.Y(_3756_), .A(regs_18__26_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf73_), );
  NAND2X1 NAND2X1_628 (.Y(_3757_), .A(_2415__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_3756_), );
  OAI21X1 OAI21X1_1491 (.Y(_3758_), .A(_3757_), .gnd(gnd), .vdd(vdd), .B(_3755_), .C(raddr1_2_bF_buf4_), );
  OAI21X1 OAI21X1_1492 (.Y(_3759_), .A(_1460_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf72_), .C(raddr1_1_bF_buf3_), );
  AOI21X1 AOI21X1_225 (.Y(_3760_), .A(regs_20__26_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf71_), .C(_3759_), );
  AND2X2 AND2X2_36 (.Y(_3761_), .A(regs_22__26_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf70_), );
  OAI21X1 OAI21X1_1493 (.Y(_3762_), .A(_1362_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf69_), .C(_2415__bF_buf3), );
  OAI21X1 OAI21X1_1494 (.Y(_3763_), .A(_3762_), .gnd(gnd), .vdd(vdd), .B(_3761_), .C(_2399__bF_buf8), );
  OAI22X1 OAI22X1_44 (.Y(_3764_), .A(_3754_), .gnd(gnd), .vdd(vdd), .B(_3758_), .C(_3763_), .D(_3760_), );
  INVX1 INVX1_135 (.Y(_3765_), .A(regs_29__26_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_629 (.Y(_3766_), .A(regs_28__26_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf68_), );
  OAI21X1 OAI21X1_1495 (.Y(_3767_), .A(_3765_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf67_), .C(_3766_), );
  MUX2X1 MUX2X1_251 (.Y(_3768_), .A(_3767_), .gnd(gnd), .vdd(vdd), .B(regs_30__26_), .S(raddr1_1_bF_buf2_), );
  NAND2X1 NAND2X1_630 (.Y(_3769_), .A(regs_26__26_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf66_), );
  OAI21X1 OAI21X1_1496 (.Y(_3770_), .A(_1195_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf65_), .C(_3769_), );
  INVX1 INVX1_136 (.Y(_3771_), .A(regs_25__26_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_631 (.Y(_3772_), .A(regs_24__26_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf64_), );
  OAI21X1 OAI21X1_1497 (.Y(_3773_), .A(_3771_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf63_), .C(_3772_), );
  MUX2X1 MUX2X1_252 (.Y(_3774_), .A(_3773_), .gnd(gnd), .vdd(vdd), .B(_3770_), .S(raddr1_1_bF_buf1_), );
  MUX2X1 MUX2X1_253 (.Y(_3775_), .A(_3774_), .gnd(gnd), .vdd(vdd), .B(_3768_), .S(raddr1_2_bF_buf3_), );
  MUX2X1 MUX2X1_254 (.Y(_3776_), .A(_3775_), .gnd(gnd), .vdd(vdd), .B(_3764_), .S(_2398__bF_buf1), );
  MUX2X1 MUX2X1_255 (.Y(_5511__26_), .A(_3752_), .gnd(gnd), .vdd(vdd), .B(_3776_), .S(raddr1_4_bF_buf3_), );
  NAND2X1 NAND2X1_632 (.Y(_3777_), .A(regs_22__27_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf62_), );
  OAI21X1 OAI21X1_1498 (.Y(_3778_), .A(_1364_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf61_), .C(_3777_), );
  NAND2X1 NAND2X1_633 (.Y(_3779_), .A(regs_20__27_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf60_), );
  OAI21X1 OAI21X1_1499 (.Y(_3780_), .A(_1462_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf59_), .C(_3779_), );
  MUX2X1 MUX2X1_256 (.Y(_3781_), .A(_3780_), .gnd(gnd), .vdd(vdd), .B(_3778_), .S(raddr1_1_bF_buf0_), );
  NAND2X1 NAND2X1_634 (.Y(_3782_), .A(_2399__bF_buf7), .gnd(gnd), .vdd(vdd), .B(_3781_), );
  NAND2X1 NAND2X1_635 (.Y(_3783_), .A(regs_18__27_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf58_), );
  OAI21X1 OAI21X1_1500 (.Y(_3784_), .A(_1561_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf57_), .C(_3783_), );
  NAND2X1 NAND2X1_636 (.Y(_3785_), .A(regs_16__27_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf56_), );
  OAI21X1 OAI21X1_1501 (.Y(_3786_), .A(_1659_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf55_), .C(_3785_), );
  MUX2X1 MUX2X1_257 (.Y(_3787_), .A(_3786_), .gnd(gnd), .vdd(vdd), .B(_3784_), .S(raddr1_1_bF_buf14_bF_buf1_), );
  AOI21X1 AOI21X1_226 (.Y(_3788_), .A(raddr1_2_bF_buf2_), .gnd(gnd), .vdd(vdd), .B(_3787_), .C(_2398__bF_buf0), );
  OAI21X1 OAI21X1_1502 (.Y(_3789_), .A(_1197_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf54_), .C(raddr1_2_bF_buf1_), );
  AOI21X1 AOI21X1_227 (.Y(_3790_), .A(regs_26__27_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf53_), .C(_3789_), );
  OAI21X1 OAI21X1_1503 (.Y(_3791_), .A(regs_30__27_), .gnd(gnd), .vdd(vdd), .B(raddr1_2_bF_buf0_), .C(_2415__bF_buf2), );
  INVX1 INVX1_137 (.Y(_3792_), .A(regs_25__27_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1504 (.Y(_3793_), .A(_3792_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf52_), .C(raddr1_2_bF_buf10_), );
  AOI21X1 AOI21X1_228 (.Y(_3794_), .A(regs_24__27_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf51_), .C(_3793_), );
  INVX1 INVX1_138 (.Y(_3795_), .A(regs_29__27_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_187 (.Y(_3796_), .A(raddr1_0_bF_buf50_), .gnd(gnd), .vdd(vdd), .B(_3795_), );
  NAND2X1 NAND2X1_637 (.Y(_3797_), .A(regs_28__27_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf49_), );
  NAND2X1 NAND2X1_638 (.Y(_3798_), .A(_2399__bF_buf6), .gnd(gnd), .vdd(vdd), .B(_3797_), );
  OAI21X1 OAI21X1_1505 (.Y(_3799_), .A(_3798_), .gnd(gnd), .vdd(vdd), .B(_3796_), .C(raddr1_1_bF_buf13_bF_buf1_), );
  OAI22X1 OAI22X1_45 (.Y(_3800_), .A(_3790_), .gnd(gnd), .vdd(vdd), .B(_3791_), .C(_3799_), .D(_3794_), );
  AOI22X1 AOI22X1_10 (.Y(_3801_), .A(_3800_), .gnd(gnd), .vdd(vdd), .B(_2398__bF_buf7), .C(_3782_), .D(_3788_), );
  NAND2X1 NAND2X1_639 (.Y(_3802_), .A(regs_6__27_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf48_), );
  OAI21X1 OAI21X1_1506 (.Y(_3803_), .A(_2155_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf47_), .C(_3802_), );
  INVX1 INVX1_139 (.Y(_3804_), .A(regs_5__27_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_640 (.Y(_3805_), .A(regs_4__27_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf46_), );
  OAI21X1 OAI21X1_1507 (.Y(_3806_), .A(_3804_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf45_), .C(_3805_), );
  MUX2X1 MUX2X1_258 (.Y(_3807_), .A(_3806_), .gnd(gnd), .vdd(vdd), .B(_3803_), .S(raddr1_1_bF_buf12_bF_buf1_), );
  INVX1 INVX1_140 (.Y(_3808_), .A(regs_3__27_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_641 (.Y(_3809_), .A(regs_2__27_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf44_), );
  OAI21X1 OAI21X1_1508 (.Y(_3810_), .A(_3808_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf43_), .C(_3809_), );
  INVX1 INVX1_141 (.Y(_3811_), .A(regs_1__27_), .gnd(gnd), .vdd(vdd), );
  NAND2X1 NAND2X1_642 (.Y(_3812_), .A(regs_0__27_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf42_), );
  OAI21X1 OAI21X1_1509 (.Y(_3813_), .A(_3811_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf41_), .C(_3812_), );
  MUX2X1 MUX2X1_259 (.Y(_3814_), .A(_3813_), .gnd(gnd), .vdd(vdd), .B(_3810_), .S(raddr1_1_bF_buf11_bF_buf1_), );
  MUX2X1 MUX2X1_260 (.Y(_3815_), .A(_3814_), .gnd(gnd), .vdd(vdd), .B(_3807_), .S(raddr1_2_bF_buf9_), );
  NAND2X1 NAND2X1_643 (.Y(_3816_), .A(regs_14__27_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf40_), );
  OAI21X1 OAI21X1_1510 (.Y(_3817_), .A(_1759_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf39_), .C(_3816_), );
  NAND2X1 NAND2X1_644 (.Y(_3818_), .A(regs_12__27_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf38_), );
  OAI21X1 OAI21X1_1511 (.Y(_3819_), .A(_1857_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf37_), .C(_3818_), );
  MUX2X1 MUX2X1_261 (.Y(_3820_), .A(_3819_), .gnd(gnd), .vdd(vdd), .B(_3817_), .S(raddr1_1_bF_buf10_bF_buf1_), );
  NAND2X1 NAND2X1_645 (.Y(_3821_), .A(regs_10__27_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf36_), );
  OAI21X1 OAI21X1_1512 (.Y(_3822_), .A(_1956_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf35_), .C(_3821_), );
  NAND2X1 NAND2X1_646 (.Y(_3823_), .A(regs_8__27_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf34_), );
  OAI21X1 OAI21X1_1513 (.Y(_3824_), .A(_2054_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf33_), .C(_3823_), );
  MUX2X1 MUX2X1_262 (.Y(_3825_), .A(_3824_), .gnd(gnd), .vdd(vdd), .B(_3822_), .S(raddr1_1_bF_buf9_bF_buf1_), );
  MUX2X1 MUX2X1_263 (.Y(_3826_), .A(_3825_), .gnd(gnd), .vdd(vdd), .B(_3820_), .S(raddr1_2_bF_buf8_), );
  MUX2X1 MUX2X1_264 (.Y(_3827_), .A(_3826_), .gnd(gnd), .vdd(vdd), .B(_3815_), .S(_2398__bF_buf6), );
  MUX2X1 MUX2X1_265 (.Y(_5511__27_), .A(_3827_), .gnd(gnd), .vdd(vdd), .B(_3801_), .S(raddr1_4_bF_buf2_), );
  NAND2X1 NAND2X1_647 (.Y(_3828_), .A(regs_22__28_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf32_), );
  OAI21X1 OAI21X1_1514 (.Y(_3829_), .A(_1366_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf31_), .C(_3828_), );
  NAND2X1 NAND2X1_648 (.Y(_3830_), .A(regs_20__28_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf30_), );
  OAI21X1 OAI21X1_1515 (.Y(_3831_), .A(_1464_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf29_), .C(_3830_), );
  MUX2X1 MUX2X1_266 (.Y(_3832_), .A(_3831_), .gnd(gnd), .vdd(vdd), .B(_3829_), .S(raddr1_1_bF_buf8_), );
  NAND2X1 NAND2X1_649 (.Y(_3833_), .A(_2399__bF_buf5), .gnd(gnd), .vdd(vdd), .B(_3832_), );
  NAND2X1 NAND2X1_650 (.Y(_3834_), .A(regs_18__28_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf28_), );
  OAI21X1 OAI21X1_1516 (.Y(_3835_), .A(_1563_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf27_), .C(_3834_), );
  NAND2X1 NAND2X1_651 (.Y(_3836_), .A(regs_16__28_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf26_), );
  OAI21X1 OAI21X1_1517 (.Y(_3837_), .A(_1661_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf25_), .C(_3836_), );
  MUX2X1 MUX2X1_267 (.Y(_3838_), .A(_3837_), .gnd(gnd), .vdd(vdd), .B(_3835_), .S(raddr1_1_bF_buf7_), );
  AOI21X1 AOI21X1_229 (.Y(_3839_), .A(raddr1_2_bF_buf7_), .gnd(gnd), .vdd(vdd), .B(_3838_), .C(_2398__bF_buf5), );
  OAI21X1 OAI21X1_1518 (.Y(_3840_), .A(_1199_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf24_), .C(raddr1_2_bF_buf6_), );
  AOI21X1 AOI21X1_230 (.Y(_3841_), .A(regs_26__28_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf23_), .C(_3840_), );
  OAI21X1 OAI21X1_1519 (.Y(_3842_), .A(regs_30__28_), .gnd(gnd), .vdd(vdd), .B(raddr1_2_bF_buf5_), .C(_2415__bF_buf1), );
  INVX1 INVX1_142 (.Y(_3843_), .A(regs_25__28_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1520 (.Y(_3844_), .A(_3843_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf22_), .C(raddr1_2_bF_buf4_), );
  AOI21X1 AOI21X1_231 (.Y(_3845_), .A(regs_24__28_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf21_), .C(_3844_), );
  INVX1 INVX1_143 (.Y(_3846_), .A(regs_29__28_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_188 (.Y(_3847_), .A(raddr1_0_bF_buf20_), .gnd(gnd), .vdd(vdd), .B(_3846_), );
  NAND2X1 NAND2X1_652 (.Y(_3848_), .A(regs_28__28_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf19_), );
  NAND2X1 NAND2X1_653 (.Y(_3849_), .A(_2399__bF_buf4), .gnd(gnd), .vdd(vdd), .B(_3848_), );
  OAI21X1 OAI21X1_1521 (.Y(_3850_), .A(_3849_), .gnd(gnd), .vdd(vdd), .B(_3847_), .C(raddr1_1_bF_buf6_), );
  OAI22X1 OAI22X1_46 (.Y(_3851_), .A(_3841_), .gnd(gnd), .vdd(vdd), .B(_3842_), .C(_3850_), .D(_3845_), );
  AOI22X1 AOI22X1_11 (.Y(_3852_), .A(_3851_), .gnd(gnd), .vdd(vdd), .B(_2398__bF_buf4), .C(_3833_), .D(_3839_), );
  INVX1 INVX1_144 (.Y(_3853_), .A(regs_5__28_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1522 (.Y(_3854_), .A(_3853_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf18_), .C(raddr1_1_bF_buf5_), );
  AOI21X1 AOI21X1_232 (.Y(_3855_), .A(regs_4__28_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf17_), .C(_3854_), );
  AND2X2 AND2X2_37 (.Y(_3856_), .A(regs_6__28_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf16_), );
  OAI21X1 OAI21X1_1523 (.Y(_3857_), .A(_2157_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf15_), .C(_2415__bF_buf0), );
  OAI21X1 OAI21X1_1524 (.Y(_3858_), .A(_3857_), .gnd(gnd), .vdd(vdd), .B(_3856_), .C(_2399__bF_buf3), );
  INVX1 INVX1_145 (.Y(_3859_), .A(regs_1__28_), .gnd(gnd), .vdd(vdd), );
  OAI21X1 OAI21X1_1525 (.Y(_3860_), .A(_3859_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf14_), .C(raddr1_1_bF_buf4_), );
  AOI21X1 AOI21X1_233 (.Y(_3861_), .A(regs_0__28_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf13_), .C(_3860_), );
  INVX1 INVX1_146 (.Y(_3862_), .A(regs_3__28_), .gnd(gnd), .vdd(vdd), );
  NOR2X1 NOR2X1_189 (.Y(_3863_), .A(raddr1_0_bF_buf12_), .gnd(gnd), .vdd(vdd), .B(_3862_), );
  NAND2X1 NAND2X1_654 (.Y(_3864_), .A(regs_2__28_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf11_), );
  NAND2X1 NAND2X1_655 (.Y(_3865_), .A(_2415__bF_buf8), .gnd(gnd), .vdd(vdd), .B(_3864_), );
  OAI21X1 OAI21X1_1526 (.Y(_3866_), .A(_3865_), .gnd(gnd), .vdd(vdd), .B(_3863_), .C(raddr1_2_bF_buf3_), );
  OAI22X1 OAI22X1_47 (.Y(_3867_), .A(_3861_), .gnd(gnd), .vdd(vdd), .B(_3866_), .C(_3858_), .D(_3855_), );
  NAND2X1 NAND2X1_656 (.Y(_3868_), .A(regs_10__28_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf10_), );
  OAI21X1 OAI21X1_1527 (.Y(_3869_), .A(_1958_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf9_), .C(_3868_), );
  NAND2X1 NAND2X1_657 (.Y(_3870_), .A(regs_8__28_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf8_), );
  OAI21X1 OAI21X1_1528 (.Y(_3871_), .A(_2056_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf7_), .C(_3870_), );
  MUX2X1 MUX2X1_268 (.Y(_3872_), .A(_3871_), .gnd(gnd), .vdd(vdd), .B(_3869_), .S(raddr1_1_bF_buf3_), );
  NAND2X1 NAND2X1_658 (.Y(_3873_), .A(regs_14__28_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf6_), );
  OAI21X1 OAI21X1_1529 (.Y(_3874_), .A(_1761_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf5_), .C(_3873_), );
  NAND2X1 NAND2X1_659 (.Y(_3875_), .A(regs_12__28_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf4_), );
  OAI21X1 OAI21X1_1530 (.Y(_3876_), .A(_1859_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf3_), .C(_3875_), );
  MUX2X1 MUX2X1_269 (.Y(_3877_), .A(_3876_), .gnd(gnd), .vdd(vdd), .B(_3874_), .S(raddr1_1_bF_buf2_), );
  MUX2X1 MUX2X1_270 (.Y(_3878_), .A(_3877_), .gnd(gnd), .vdd(vdd), .B(_3872_), .S(_2399__bF_buf2), );
  MUX2X1 MUX2X1_271 (.Y(_3879_), .A(_3878_), .gnd(gnd), .vdd(vdd), .B(_3867_), .S(_2398__bF_buf3), );
  MUX2X1 MUX2X1_272 (.Y(_5511__28_), .A(_3879_), .gnd(gnd), .vdd(vdd), .B(_3852_), .S(raddr1_4_bF_buf1_), );
  NAND2X1 NAND2X1_660 (.Y(_3880_), .A(regs_22__29_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf2_), );
  OAI21X1 OAI21X1_1531 (.Y(_3881_), .A(_1368_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf1_), .C(_3880_), );
  NAND2X1 NAND2X1_661 (.Y(_3882_), .A(regs_20__29_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf0_), );
  OAI21X1 OAI21X1_1532 (.Y(_3883_), .A(_1466_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf96_), .C(_3882_), );
  MUX2X1 MUX2X1_273 (.Y(_3884_), .A(_3883_), .gnd(gnd), .vdd(vdd), .B(_3881_), .S(raddr1_1_bF_buf1_), );
  NAND2X1 NAND2X1_662 (.Y(_3885_), .A(_2399__bF_buf1), .gnd(gnd), .vdd(vdd), .B(_3884_), );
  NAND2X1 NAND2X1_663 (.Y(_3886_), .A(regs_18__29_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf95_), );
  OAI21X1 OAI21X1_1533 (.Y(_3887_), .A(_1565_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf94_), .C(_3886_), );
  NAND2X1 NAND2X1_664 (.Y(_3888_), .A(regs_16__29_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf93_), );
  OAI21X1 OAI21X1_1534 (.Y(_3889_), .A(_1663_), .gnd(gnd), .vdd(vdd), .B(raddr1_0_bF_buf92_), .C(_3888_), );
  MUX2X1 MUX2X1_274 (.gnd(gnd), .A(_3889_), .Y(_3890_), .vdd(vdd), .B(_3887_), .S(raddr1_1_bF_buf0_), );
  AOI21X1 AOI21X1_234 (.gnd(gnd), .A(raddr1_2_bF_buf2_), .Y(_3891_), .vdd(vdd), .B(_3890_), .C(_2398__bF_buf2), );
  OAI21X1 OAI21X1_1535 (.gnd(gnd), .A(_1201_), .Y(_3892_), .vdd(vdd), .B(raddr1_0_bF_buf91_), .C(raddr1_2_bF_buf1_), );
  AOI21X1 AOI21X1_235 (.gnd(gnd), .A(regs_26__29_), .Y(_3893_), .vdd(vdd), .B(raddr1_0_bF_buf90_), .C(_3892_), );
  OAI21X1 OAI21X1_1536 (.gnd(gnd), .A(regs_30__29_), .Y(_3894_), .vdd(vdd), .B(raddr1_2_bF_buf0_), .C(_2415__bF_buf7), );
  INVX1 INVX1_147 (.gnd(gnd), .A(regs_25__29_), .Y(_3895_), .vdd(vdd), );
  OAI21X1 OAI21X1_1537 (.gnd(gnd), .A(_3895_), .Y(_3896_), .vdd(vdd), .B(raddr1_0_bF_buf89_), .C(raddr1_2_bF_buf10_), );
  AOI21X1 AOI21X1_236 (.gnd(gnd), .A(regs_24__29_), .Y(_3897_), .vdd(vdd), .B(raddr1_0_bF_buf88_), .C(_3896_), );
  INVX1 INVX1_148 (.gnd(gnd), .A(regs_29__29_), .Y(_3898_), .vdd(vdd), );
  NOR2X1 NOR2X1_190 (.gnd(gnd), .A(raddr1_0_bF_buf87_), .Y(_3899_), .vdd(vdd), .B(_3898_), );
  NAND2X1 NAND2X1_665 (.gnd(gnd), .A(regs_28__29_), .Y(_3900_), .vdd(vdd), .B(raddr1_0_bF_buf86_), );
  NAND2X1 NAND2X1_666 (.gnd(gnd), .A(_2399__bF_buf0), .Y(_3901_), .vdd(vdd), .B(_3900_), );
  OAI21X1 OAI21X1_1538 (.gnd(gnd), .A(_3901_), .Y(_3902_), .vdd(vdd), .B(_3899_), .C(raddr1_1_bF_buf14_bF_buf0_), );
  OAI22X1 OAI22X1_48 (.gnd(gnd), .A(_3893_), .Y(_3903_), .vdd(vdd), .B(_3894_), .C(_3902_), .D(_3897_), );
  AOI22X1 AOI22X1_12 (.gnd(gnd), .A(_3903_), .Y(_3904_), .vdd(vdd), .B(_2398__bF_buf1), .C(_3885_), .D(_3891_), );
  INVX1 INVX1_149 (.gnd(gnd), .A(regs_5__29_), .Y(_3905_), .vdd(vdd), );
  OAI21X1 OAI21X1_1539 (.gnd(gnd), .A(_3905_), .Y(_3906_), .vdd(vdd), .B(raddr1_0_bF_buf85_), .C(raddr1_1_bF_buf13_bF_buf0_), );
  AOI21X1 AOI21X1_237 (.gnd(gnd), .A(regs_4__29_), .Y(_3907_), .vdd(vdd), .B(raddr1_0_bF_buf84_), .C(_3906_), );
  AND2X2 AND2X2_38 (.gnd(gnd), .A(regs_6__29_), .Y(_3908_), .vdd(vdd), .B(raddr1_0_bF_buf83_), );
  OAI21X1 OAI21X1_1540 (.gnd(gnd), .A(_2159_), .Y(_3909_), .vdd(vdd), .B(raddr1_0_bF_buf82_), .C(_2415__bF_buf6), );
  OAI21X1 OAI21X1_1541 (.gnd(gnd), .A(_3909_), .Y(_3910_), .vdd(vdd), .B(_3908_), .C(_2399__bF_buf8), );
  INVX1 INVX1_150 (.gnd(gnd), .A(regs_1__29_), .Y(_3911_), .vdd(vdd), );
  OAI21X1 OAI21X1_1542 (.gnd(gnd), .A(_3911_), .Y(_3912_), .vdd(vdd), .B(raddr1_0_bF_buf81_), .C(raddr1_1_bF_buf12_bF_buf0_), );
  AOI21X1 AOI21X1_238 (.gnd(gnd), .A(regs_0__29_), .Y(_3913_), .vdd(vdd), .B(raddr1_0_bF_buf80_), .C(_3912_), );
  INVX1 INVX1_151 (.gnd(gnd), .A(regs_3__29_), .Y(_3914_), .vdd(vdd), );
  NOR2X1 NOR2X1_191 (.gnd(gnd), .A(raddr1_0_bF_buf79_), .Y(_3915_), .vdd(vdd), .B(_3914_), );
  NAND2X1 NAND2X1_667 (.gnd(gnd), .A(regs_2__29_), .Y(_3916_), .vdd(vdd), .B(raddr1_0_bF_buf78_), );
  NAND2X1 NAND2X1_668 (.gnd(gnd), .A(_2415__bF_buf5), .Y(_3917_), .vdd(vdd), .B(_3916_), );
  OAI21X1 OAI21X1_1543 (.gnd(gnd), .A(_3917_), .Y(_3918_), .vdd(vdd), .B(_3915_), .C(raddr1_2_bF_buf9_), );
  OAI22X1 OAI22X1_49 (.gnd(gnd), .A(_3913_), .Y(_3919_), .vdd(vdd), .B(_3918_), .C(_3910_), .D(_3907_), );
  NAND2X1 NAND2X1_669 (.gnd(gnd), .A(regs_10__29_), .Y(_3920_), .vdd(vdd), .B(raddr1_0_bF_buf77_), );
  OAI21X1 OAI21X1_1544 (.gnd(gnd), .A(_1960_), .Y(_3921_), .vdd(vdd), .B(raddr1_0_bF_buf76_), .C(_3920_), );
  NAND2X1 NAND2X1_670 (.gnd(gnd), .A(regs_8__29_), .Y(_3922_), .vdd(vdd), .B(raddr1_0_bF_buf75_), );
  OAI21X1 OAI21X1_1545 (.gnd(gnd), .A(_2058_), .Y(_3923_), .vdd(vdd), .B(raddr1_0_bF_buf74_), .C(_3922_), );
  MUX2X1 MUX2X1_275 (.gnd(gnd), .A(_3923_), .Y(_3924_), .vdd(vdd), .B(_3921_), .S(raddr1_1_bF_buf11_bF_buf0_), );
  NAND2X1 NAND2X1_671 (.gnd(gnd), .A(regs_14__29_), .Y(_3925_), .vdd(vdd), .B(raddr1_0_bF_buf73_), );
  OAI21X1 OAI21X1_1546 (.gnd(gnd), .A(_1763_), .Y(_3926_), .vdd(vdd), .B(raddr1_0_bF_buf72_), .C(_3925_), );
  NAND2X1 NAND2X1_672 (.gnd(gnd), .A(regs_12__29_), .Y(_3927_), .vdd(vdd), .B(raddr1_0_bF_buf71_), );
  OAI21X1 OAI21X1_1547 (.gnd(gnd), .A(_1861_), .Y(_3928_), .vdd(vdd), .B(raddr1_0_bF_buf70_), .C(_3927_), );
  MUX2X1 MUX2X1_276 (.gnd(gnd), .A(_3928_), .Y(_3929_), .vdd(vdd), .B(_3926_), .S(raddr1_1_bF_buf10_bF_buf0_), );
  MUX2X1 MUX2X1_277 (.gnd(gnd), .A(_3929_), .Y(_3930_), .vdd(vdd), .B(_3924_), .S(_2399__bF_buf7), );
  MUX2X1 MUX2X1_278 (.gnd(gnd), .A(_3930_), .Y(_3931_), .vdd(vdd), .B(_3919_), .S(_2398__bF_buf0), );
  MUX2X1 MUX2X1_279 (.gnd(gnd), .A(_3931_), .Y(_5511__29_), .vdd(vdd), .B(_3904_), .S(raddr1_4_bF_buf0_), );
  OAI21X1 OAI21X1_1548 (.gnd(gnd), .A(_1468_), .Y(_3932_), .vdd(vdd), .B(raddr1_0_bF_buf69_), .C(raddr1_1_bF_buf9_bF_buf0_), );
  AOI21X1 AOI21X1_239 (.gnd(gnd), .A(regs_20__30_), .Y(_3933_), .vdd(vdd), .B(raddr1_0_bF_buf68_), .C(_3932_), );
  AND2X2 AND2X2_39 (.gnd(gnd), .A(regs_22__30_), .Y(_3934_), .vdd(vdd), .B(raddr1_0_bF_buf67_), );
  OAI21X1 OAI21X1_1549 (.gnd(gnd), .A(_1370_), .Y(_3935_), .vdd(vdd), .B(raddr1_0_bF_buf66_), .C(_2415__bF_buf4), );
  OAI21X1 OAI21X1_1550 (.gnd(gnd), .A(_3935_), .Y(_3936_), .vdd(vdd), .B(_3934_), .C(_2399__bF_buf6), );
  OAI21X1 OAI21X1_1551 (.gnd(gnd), .A(_1665_), .Y(_3937_), .vdd(vdd), .B(raddr1_0_bF_buf65_), .C(raddr1_1_bF_buf8_), );
  AOI21X1 AOI21X1_240 (.gnd(gnd), .A(regs_16__30_), .Y(_3938_), .vdd(vdd), .B(raddr1_0_bF_buf64_), .C(_3937_), );
  NOR2X1 NOR2X1_192 (.gnd(gnd), .A(raddr1_0_bF_buf63_), .Y(_3939_), .vdd(vdd), .B(_1567_), );
  NAND2X1 NAND2X1_673 (.gnd(gnd), .A(regs_18__30_), .Y(_3940_), .vdd(vdd), .B(raddr1_0_bF_buf62_), );
  NAND2X1 NAND2X1_674 (.gnd(gnd), .A(_2415__bF_buf3), .Y(_3941_), .vdd(vdd), .B(_3940_), );
  OAI21X1 OAI21X1_1552 (.gnd(gnd), .A(_3941_), .Y(_3942_), .vdd(vdd), .B(_3939_), .C(raddr1_2_bF_buf8_), );
  OAI22X1 OAI22X1_50 (.gnd(gnd), .A(_3938_), .Y(_3943_), .vdd(vdd), .B(_3942_), .C(_3936_), .D(_3933_), );
  INVX1 INVX1_152 (.gnd(gnd), .A(regs_29__30_), .Y(_3944_), .vdd(vdd), );
  NAND2X1 NAND2X1_675 (.gnd(gnd), .A(regs_28__30_), .Y(_3945_), .vdd(vdd), .B(raddr1_0_bF_buf61_), );
  OAI21X1 OAI21X1_1553 (.gnd(gnd), .A(_3944_), .Y(_3946_), .vdd(vdd), .B(raddr1_0_bF_buf60_), .C(_3945_), );
  MUX2X1 MUX2X1_280 (.gnd(gnd), .A(_3946_), .Y(_3947_), .vdd(vdd), .B(regs_30__30_), .S(raddr1_1_bF_buf7_), );
  NAND2X1 NAND2X1_676 (.gnd(gnd), .A(regs_26__30_), .Y(_3948_), .vdd(vdd), .B(raddr1_0_bF_buf59_), );
  OAI21X1 OAI21X1_1554 (.gnd(gnd), .A(_1203_), .Y(_3949_), .vdd(vdd), .B(raddr1_0_bF_buf58_), .C(_3948_), );
  INVX1 INVX1_153 (.gnd(gnd), .A(regs_25__30_), .Y(_3950_), .vdd(vdd), );
  NAND2X1 NAND2X1_677 (.gnd(gnd), .A(regs_24__30_), .Y(_3951_), .vdd(vdd), .B(raddr1_0_bF_buf57_), );
  OAI21X1 OAI21X1_1555 (.gnd(gnd), .A(_3950_), .Y(_3952_), .vdd(vdd), .B(raddr1_0_bF_buf56_), .C(_3951_), );
  MUX2X1 MUX2X1_281 (.gnd(gnd), .A(_3952_), .Y(_3953_), .vdd(vdd), .B(_3949_), .S(raddr1_1_bF_buf6_), );
  MUX2X1 MUX2X1_282 (.gnd(gnd), .A(_3953_), .Y(_3954_), .vdd(vdd), .B(_3947_), .S(raddr1_2_bF_buf7_), );
  MUX2X1 MUX2X1_283 (.gnd(gnd), .A(_3954_), .Y(_3955_), .vdd(vdd), .B(_3943_), .S(_2398__bF_buf7), );
  NAND2X1 NAND2X1_678 (.gnd(gnd), .A(regs_6__30_), .Y(_3956_), .vdd(vdd), .B(raddr1_0_bF_buf55_), );
  OAI21X1 OAI21X1_1556 (.gnd(gnd), .A(_2161_), .Y(_3957_), .vdd(vdd), .B(raddr1_0_bF_buf54_), .C(_3956_), );
  INVX1 INVX1_154 (.gnd(gnd), .A(regs_5__30_), .Y(_3958_), .vdd(vdd), );
  NAND2X1 NAND2X1_679 (.gnd(gnd), .A(regs_4__30_), .Y(_3959_), .vdd(vdd), .B(raddr1_0_bF_buf53_), );
  OAI21X1 OAI21X1_1557 (.gnd(gnd), .A(_3958_), .Y(_3960_), .vdd(vdd), .B(raddr1_0_bF_buf52_), .C(_3959_), );
  MUX2X1 MUX2X1_284 (.gnd(gnd), .A(_3960_), .Y(_3961_), .vdd(vdd), .B(_3957_), .S(raddr1_1_bF_buf5_), );
  INVX1 INVX1_155 (.gnd(gnd), .A(regs_3__30_), .Y(_3962_), .vdd(vdd), );
  NAND2X1 NAND2X1_680 (.gnd(gnd), .A(regs_2__30_), .Y(_3963_), .vdd(vdd), .B(raddr1_0_bF_buf51_), );
  OAI21X1 OAI21X1_1558 (.gnd(gnd), .A(_3962_), .Y(_3964_), .vdd(vdd), .B(raddr1_0_bF_buf50_), .C(_3963_), );
  INVX1 INVX1_156 (.gnd(gnd), .A(regs_1__30_), .Y(_3965_), .vdd(vdd), );
  NAND2X1 NAND2X1_681 (.gnd(gnd), .A(regs_0__30_), .Y(_3966_), .vdd(vdd), .B(raddr1_0_bF_buf49_), );
  OAI21X1 OAI21X1_1559 (.gnd(gnd), .A(_3965_), .Y(_3967_), .vdd(vdd), .B(raddr1_0_bF_buf48_), .C(_3966_), );
  MUX2X1 MUX2X1_285 (.gnd(gnd), .A(_3967_), .Y(_3968_), .vdd(vdd), .B(_3964_), .S(raddr1_1_bF_buf4_), );
  MUX2X1 MUX2X1_286 (.gnd(gnd), .A(_3968_), .Y(_3969_), .vdd(vdd), .B(_3961_), .S(raddr1_2_bF_buf6_), );
  NAND2X1 NAND2X1_682 (.gnd(gnd), .A(regs_10__30_), .Y(_3970_), .vdd(vdd), .B(raddr1_0_bF_buf47_), );
  OAI21X1 OAI21X1_1560 (.gnd(gnd), .A(_1962_), .Y(_3971_), .vdd(vdd), .B(raddr1_0_bF_buf46_), .C(_3970_), );
  NAND2X1 NAND2X1_683 (.gnd(gnd), .A(regs_8__30_), .Y(_3972_), .vdd(vdd), .B(raddr1_0_bF_buf45_), );
  OAI21X1 OAI21X1_1561 (.gnd(gnd), .A(_2060_), .Y(_3973_), .vdd(vdd), .B(raddr1_0_bF_buf44_), .C(_3972_), );
  MUX2X1 MUX2X1_287 (.gnd(gnd), .A(_3973_), .Y(_3974_), .vdd(vdd), .B(_3971_), .S(raddr1_1_bF_buf3_), );
  NAND2X1 NAND2X1_684 (.gnd(gnd), .A(regs_14__30_), .Y(_3975_), .vdd(vdd), .B(raddr1_0_bF_buf43_), );
  OAI21X1 OAI21X1_1562 (.gnd(gnd), .A(_1765_), .Y(_3976_), .vdd(vdd), .B(raddr1_0_bF_buf42_), .C(_3975_), );
  NAND2X1 NAND2X1_685 (.gnd(gnd), .A(regs_12__30_), .Y(_3977_), .vdd(vdd), .B(raddr1_0_bF_buf41_), );
  OAI21X1 OAI21X1_1563 (.gnd(gnd), .A(_1863_), .Y(_3978_), .vdd(vdd), .B(raddr1_0_bF_buf40_), .C(_3977_), );
  MUX2X1 MUX2X1_288 (.gnd(gnd), .A(_3978_), .Y(_3979_), .vdd(vdd), .B(_3976_), .S(raddr1_1_bF_buf2_), );
  MUX2X1 MUX2X1_289 (.gnd(gnd), .A(_3979_), .Y(_3980_), .vdd(vdd), .B(_3974_), .S(_2399__bF_buf5), );
  MUX2X1 MUX2X1_290 (.gnd(gnd), .A(_3980_), .Y(_3981_), .vdd(vdd), .B(_3969_), .S(_2398__bF_buf6), );
  MUX2X1 MUX2X1_291 (.gnd(gnd), .A(_3981_), .Y(_5511__30_), .vdd(vdd), .B(_3955_), .S(raddr1_4_bF_buf4_), );
  INVX1 INVX1_157 (.gnd(gnd), .A(regs_5__31_), .Y(_3982_), .vdd(vdd), );
  OAI21X1 OAI21X1_1564 (.gnd(gnd), .A(_3982_), .Y(_3983_), .vdd(vdd), .B(raddr1_0_bF_buf39_), .C(raddr1_1_bF_buf1_), );
  AOI21X1 AOI21X1_241 (.gnd(gnd), .A(regs_4__31_), .Y(_3984_), .vdd(vdd), .B(raddr1_0_bF_buf38_), .C(_3983_), );
  AND2X2 AND2X2_40 (.gnd(gnd), .A(regs_6__31_), .Y(_3985_), .vdd(vdd), .B(raddr1_0_bF_buf37_), );
  OAI21X1 OAI21X1_1565 (.gnd(gnd), .A(_2163_), .Y(_3986_), .vdd(vdd), .B(raddr1_0_bF_buf36_), .C(_2415__bF_buf2), );
  OAI21X1 OAI21X1_1566 (.gnd(gnd), .A(_3986_), .Y(_3987_), .vdd(vdd), .B(_3985_), .C(_2399__bF_buf4), );
  INVX1 INVX1_158 (.gnd(gnd), .A(regs_1__31_), .Y(_3988_), .vdd(vdd), );
  OAI21X1 OAI21X1_1567 (.gnd(gnd), .A(_3988_), .Y(_3989_), .vdd(vdd), .B(raddr1_0_bF_buf35_), .C(raddr1_1_bF_buf0_), );
  AOI21X1 AOI21X1_242 (.gnd(gnd), .A(regs_0__31_), .Y(_3990_), .vdd(vdd), .B(raddr1_0_bF_buf34_), .C(_3989_), );
  INVX1 INVX1_159 (.gnd(gnd), .A(regs_3__31_), .Y(_3991_), .vdd(vdd), );
  NOR2X1 NOR2X1_193 (.gnd(gnd), .A(raddr1_0_bF_buf33_), .Y(_3992_), .vdd(vdd), .B(_3991_), );
  NAND2X1 NAND2X1_686 (.gnd(gnd), .A(regs_2__31_), .Y(_3993_), .vdd(vdd), .B(raddr1_0_bF_buf32_), );
  NAND2X1 NAND2X1_687 (.gnd(gnd), .A(_2415__bF_buf1), .Y(_3994_), .vdd(vdd), .B(_3993_), );
  OAI21X1 OAI21X1_1568 (.gnd(gnd), .A(_3994_), .Y(_3995_), .vdd(vdd), .B(_3992_), .C(raddr1_2_bF_buf5_), );
  OAI22X1 OAI22X1_51 (.gnd(gnd), .A(_3990_), .Y(_3996_), .vdd(vdd), .B(_3995_), .C(_3987_), .D(_3984_), );
  NAND2X1 NAND2X1_688 (.gnd(gnd), .A(regs_10__31_), .Y(_3997_), .vdd(vdd), .B(raddr1_0_bF_buf31_), );
  OAI21X1 OAI21X1_1569 (.gnd(gnd), .A(_1964_), .Y(_3998_), .vdd(vdd), .B(raddr1_0_bF_buf30_), .C(_3997_), );
  NAND2X1 NAND2X1_689 (.gnd(gnd), .A(regs_8__31_), .Y(_3999_), .vdd(vdd), .B(raddr1_0_bF_buf29_), );
  OAI21X1 OAI21X1_1570 (.gnd(gnd), .A(_2062_), .Y(_4000_), .vdd(vdd), .B(raddr1_0_bF_buf28_), .C(_3999_), );
  MUX2X1 MUX2X1_292 (.gnd(gnd), .A(_4000_), .Y(_4001_), .vdd(vdd), .B(_3998_), .S(raddr1_1_bF_buf14_bF_buf3_), );
  NAND2X1 NAND2X1_690 (.gnd(gnd), .A(regs_14__31_), .Y(_4002_), .vdd(vdd), .B(raddr1_0_bF_buf27_), );
  OAI21X1 OAI21X1_1571 (.gnd(gnd), .A(_1767_), .Y(_4003_), .vdd(vdd), .B(raddr1_0_bF_buf26_), .C(_4002_), );
  NAND2X1 NAND2X1_691 (.gnd(gnd), .A(regs_12__31_), .Y(_4004_), .vdd(vdd), .B(raddr1_0_bF_buf25_), );
  OAI21X1 OAI21X1_1572 (.gnd(gnd), .A(_1865_), .Y(_4005_), .vdd(vdd), .B(raddr1_0_bF_buf24_), .C(_4004_), );
  MUX2X1 MUX2X1_293 (.gnd(gnd), .A(_4005_), .Y(_4006_), .vdd(vdd), .B(_4003_), .S(raddr1_1_bF_buf13_bF_buf3_), );
  MUX2X1 MUX2X1_294 (.gnd(gnd), .A(_4006_), .Y(_4007_), .vdd(vdd), .B(_4001_), .S(_2399__bF_buf3), );
  MUX2X1 MUX2X1_295 (.gnd(gnd), .A(_4007_), .Y(_4008_), .vdd(vdd), .B(_3996_), .S(_2398__bF_buf5), );
  OAI21X1 OAI21X1_1573 (.gnd(gnd), .A(_1667_), .Y(_4009_), .vdd(vdd), .B(raddr1_0_bF_buf23_), .C(raddr1_1_bF_buf12_bF_buf3_), );
  AOI21X1 AOI21X1_243 (.gnd(gnd), .A(regs_16__31_), .Y(_4010_), .vdd(vdd), .B(raddr1_0_bF_buf22_), .C(_4009_), );
  NOR2X1 NOR2X1_194 (.gnd(gnd), .A(raddr1_0_bF_buf21_), .Y(_4011_), .vdd(vdd), .B(_1569_), );
  NAND2X1 NAND2X1_692 (.gnd(gnd), .A(regs_18__31_), .Y(_4012_), .vdd(vdd), .B(raddr1_0_bF_buf20_), );
  NAND2X1 NAND2X1_693 (.gnd(gnd), .A(_2415__bF_buf0), .Y(_4013_), .vdd(vdd), .B(_4012_), );
  OAI21X1 OAI21X1_1574 (.gnd(gnd), .A(_4013_), .Y(_4014_), .vdd(vdd), .B(_4011_), .C(raddr1_2_bF_buf4_), );
  OAI21X1 OAI21X1_1575 (.gnd(gnd), .A(_1470_), .Y(_4015_), .vdd(vdd), .B(raddr1_0_bF_buf19_), .C(raddr1_1_bF_buf11_bF_buf3_), );
  AOI21X1 AOI21X1_244 (.gnd(gnd), .A(regs_20__31_), .Y(_4016_), .vdd(vdd), .B(raddr1_0_bF_buf18_), .C(_4015_), );
  AND2X2 AND2X2_41 (.gnd(gnd), .A(regs_22__31_), .Y(_4017_), .vdd(vdd), .B(raddr1_0_bF_buf17_), );
  OAI21X1 OAI21X1_1576 (.gnd(gnd), .A(_1372_), .Y(_4018_), .vdd(vdd), .B(raddr1_0_bF_buf16_), .C(_2415__bF_buf8), );
  OAI21X1 OAI21X1_1577 (.gnd(gnd), .A(_4018_), .Y(_4019_), .vdd(vdd), .B(_4017_), .C(_2399__bF_buf2), );
  OAI22X1 OAI22X1_52 (.gnd(gnd), .A(_4010_), .Y(_4020_), .vdd(vdd), .B(_4014_), .C(_4019_), .D(_4016_), );
  INVX1 INVX1_160 (.gnd(gnd), .A(regs_29__31_), .Y(_4021_), .vdd(vdd), );
  NAND2X1 NAND2X1_694 (.gnd(gnd), .A(regs_28__31_), .Y(_4022_), .vdd(vdd), .B(raddr1_0_bF_buf15_), );
  OAI21X1 OAI21X1_1578 (.gnd(gnd), .A(_4021_), .Y(_4023_), .vdd(vdd), .B(raddr1_0_bF_buf14_), .C(_4022_), );
  MUX2X1 MUX2X1_296 (.gnd(gnd), .A(_4023_), .Y(_4024_), .vdd(vdd), .B(regs_30__31_), .S(raddr1_1_bF_buf10_bF_buf3_), );
  NAND2X1 NAND2X1_695 (.gnd(gnd), .A(regs_26__31_), .Y(_4025_), .vdd(vdd), .B(raddr1_0_bF_buf13_), );
  OAI21X1 OAI21X1_1579 (.gnd(gnd), .A(_1205_), .Y(_4026_), .vdd(vdd), .B(raddr1_0_bF_buf12_), .C(_4025_), );
  INVX1 INVX1_161 (.gnd(gnd), .A(regs_25__31_), .Y(_4027_), .vdd(vdd), );
  NAND2X1 NAND2X1_696 (.gnd(gnd), .A(regs_24__31_), .Y(_4028_), .vdd(vdd), .B(raddr1_0_bF_buf11_), );
  OAI21X1 OAI21X1_1580 (.gnd(gnd), .A(_4027_), .Y(_4029_), .vdd(vdd), .B(raddr1_0_bF_buf10_), .C(_4028_), );
  MUX2X1 MUX2X1_297 (.gnd(gnd), .A(_4029_), .Y(_4030_), .vdd(vdd), .B(_4026_), .S(raddr1_1_bF_buf9_bF_buf3_), );
  MUX2X1 MUX2X1_298 (.gnd(gnd), .A(_4030_), .Y(_4031_), .vdd(vdd), .B(_4024_), .S(raddr1_2_bF_buf3_), );
  MUX2X1 MUX2X1_299 (.gnd(gnd), .A(_4031_), .Y(_4032_), .vdd(vdd), .B(_4020_), .S(_2398__bF_buf4), );
  MUX2X1 MUX2X1_300 (.gnd(gnd), .A(_4008_), .Y(_5511__31_), .vdd(vdd), .B(_4032_), .S(raddr1_4_bF_buf3_), );
  INVX8 INVX8_5 (.gnd(gnd), .A(raddr2[3]), .Y(_4033_), .vdd(vdd), );
  OAI21X1 OAI21X1_1581 (.gnd(gnd), .A(_2427_), .Y(_4034_), .vdd(vdd), .B(raddr2_0_bF_buf96_), .C(raddr2_1_bF_buf14_bF_buf3_), );
  AOI21X1 AOI21X1_245 (.gnd(gnd), .A(regs_4__0_), .Y(_4035_), .vdd(vdd), .B(raddr2_0_bF_buf95_), .C(_4034_), );
  INVX8 INVX8_6 (.gnd(gnd), .A(raddr2_2_bF_buf10_), .Y(_4036_), .vdd(vdd), );
  AND2X2 AND2X2_42 (.gnd(gnd), .A(regs_6__0_), .Y(_4037_), .vdd(vdd), .B(raddr2_0_bF_buf94_), );
  INVX8 INVX8_7 (.gnd(gnd), .A(raddr2_1_bF_buf13_bF_buf3_), .Y(_4038_), .vdd(vdd), );
  OAI21X1 OAI21X1_1582 (.gnd(gnd), .A(_2097_), .Y(_4039_), .vdd(vdd), .B(raddr2_0_bF_buf93_), .C(_4038__bF_buf8), );
  OAI21X1 OAI21X1_1583 (.gnd(gnd), .A(_4039_), .Y(_4040_), .vdd(vdd), .B(_4037_), .C(_4036__bF_buf8), );
  OAI21X1 OAI21X1_1584 (.gnd(gnd), .A(_2433_), .Y(_4041_), .vdd(vdd), .B(raddr2_0_bF_buf92_), .C(raddr2_1_bF_buf12_bF_buf3_), );
  AOI21X1 AOI21X1_246 (.gnd(gnd), .A(regs_0__0_), .Y(_4042_), .vdd(vdd), .B(raddr2_0_bF_buf91_), .C(_4041_), );
  AOI21X1 AOI21X1_247 (.gnd(gnd), .A(regs_2__0_), .Y(_4043_), .vdd(vdd), .B(raddr2_0_bF_buf90_), .C(raddr2_1_bF_buf11_), );
  OAI21X1 OAI21X1_1585 (.gnd(gnd), .A(_2436_), .Y(_4044_), .vdd(vdd), .B(raddr2_0_bF_buf89_), .C(_4043_), );
  NAND2X1 NAND2X1_697 (.gnd(gnd), .A(raddr2_2_bF_buf9_), .Y(_4045_), .vdd(vdd), .B(_4044_), );
  OAI22X1 OAI22X1_53 (.gnd(gnd), .A(_4045_), .Y(_4046_), .vdd(vdd), .B(_4042_), .C(_4040_), .D(_4035_), );
  NAND2X1 NAND2X1_698 (.gnd(gnd), .A(regs_10__0_), .Y(_4047_), .vdd(vdd), .B(raddr2_0_bF_buf88_), );
  OAI21X1 OAI21X1_1586 (.gnd(gnd), .A(_1900_), .Y(_4048_), .vdd(vdd), .B(raddr2_0_bF_buf87_), .C(_4047_), );
  NAND2X1 NAND2X1_699 (.gnd(gnd), .A(regs_8__0_), .Y(_4049_), .vdd(vdd), .B(raddr2_0_bF_buf86_), );
  OAI21X1 OAI21X1_1587 (.gnd(gnd), .A(_1999_), .Y(_4050_), .vdd(vdd), .B(raddr2_0_bF_buf85_), .C(_4049_), );
  MUX2X1 MUX2X1_301 (.gnd(gnd), .A(_4050_), .Y(_4051_), .vdd(vdd), .B(_4048_), .S(raddr2_1_bF_buf10_), );
  NAND2X1 NAND2X1_700 (.gnd(gnd), .A(regs_14__0_), .Y(_4052_), .vdd(vdd), .B(raddr2_0_bF_buf84_), );
  OAI21X1 OAI21X1_1588 (.gnd(gnd), .A(_1702_), .Y(_4053_), .vdd(vdd), .B(raddr2_0_bF_buf83_), .C(_4052_), );
  NAND2X1 NAND2X1_701 (.gnd(gnd), .A(regs_12__0_), .Y(_4054_), .vdd(vdd), .B(raddr2_0_bF_buf82_), );
  OAI21X1 OAI21X1_1589 (.gnd(gnd), .A(_1802_), .Y(_4055_), .vdd(vdd), .B(raddr2_0_bF_buf81_), .C(_4054_), );
  MUX2X1 MUX2X1_302 (.gnd(gnd), .A(_4055_), .Y(_4056_), .vdd(vdd), .B(_4053_), .S(raddr2_1_bF_buf9_), );
  MUX2X1 MUX2X1_303 (.gnd(gnd), .A(_4056_), .Y(_4057_), .vdd(vdd), .B(_4051_), .S(_4036__bF_buf7), );
  MUX2X1 MUX2X1_304 (.gnd(gnd), .A(_4057_), .Y(_4058_), .vdd(vdd), .B(_4046_), .S(_4033__bF_buf7), );
  OAI21X1 OAI21X1_1590 (.gnd(gnd), .A(_1604_), .Y(_4059_), .vdd(vdd), .B(raddr2_0_bF_buf80_), .C(raddr2_1_bF_buf8_), );
  AOI21X1 AOI21X1_248 (.gnd(gnd), .A(regs_16__0_), .Y(_4060_), .vdd(vdd), .B(raddr2_0_bF_buf79_), .C(_4059_), );
  NOR2X1 NOR2X1_195 (.gnd(gnd), .A(raddr2_0_bF_buf78_), .Y(_4061_), .vdd(vdd), .B(_1505_), );
  NAND2X1 NAND2X1_702 (.gnd(gnd), .A(regs_18__0_), .Y(_4062_), .vdd(vdd), .B(raddr2_0_bF_buf77_), );
  NAND2X1 NAND2X1_703 (.gnd(gnd), .A(_4038__bF_buf7), .Y(_4063_), .vdd(vdd), .B(_4062_), );
  OAI21X1 OAI21X1_1591 (.gnd(gnd), .A(_4063_), .Y(_4064_), .vdd(vdd), .B(_4061_), .C(raddr2_2_bF_buf8_), );
  OAI21X1 OAI21X1_1592 (.gnd(gnd), .A(_1407_), .Y(_4065_), .vdd(vdd), .B(raddr2_0_bF_buf76_), .C(raddr2_1_bF_buf7_), );
  AOI21X1 AOI21X1_249 (.gnd(gnd), .A(regs_20__0_), .Y(_4066_), .vdd(vdd), .B(raddr2_0_bF_buf75_), .C(_4065_), );
  AND2X2 AND2X2_43 (.gnd(gnd), .A(regs_22__0_), .Y(_4067_), .vdd(vdd), .B(raddr2_0_bF_buf74_), );
  OAI21X1 OAI21X1_1593 (.gnd(gnd), .A(_1307_), .Y(_4068_), .vdd(vdd), .B(raddr2_0_bF_buf73_), .C(_4038__bF_buf6), );
  OAI21X1 OAI21X1_1594 (.gnd(gnd), .A(_4068_), .Y(_4069_), .vdd(vdd), .B(_4067_), .C(_4036__bF_buf6), );
  OAI22X1 OAI22X1_54 (.gnd(gnd), .A(_4060_), .Y(_4070_), .vdd(vdd), .B(_4064_), .C(_4069_), .D(_4066_), );
  NAND2X1 NAND2X1_704 (.gnd(gnd), .A(regs_28__0_), .Y(_4071_), .vdd(vdd), .B(raddr2_0_bF_buf72_), );
  OAI21X1 OAI21X1_1595 (.gnd(gnd), .A(_2420_), .Y(_4072_), .vdd(vdd), .B(raddr2_0_bF_buf71_), .C(_4071_), );
  MUX2X1 MUX2X1_305 (.gnd(gnd), .A(_4072_), .Y(_4073_), .vdd(vdd), .B(regs_30__0_), .S(raddr2_1_bF_buf6_), );
  NAND2X1 NAND2X1_705 (.gnd(gnd), .A(regs_26__0_), .Y(_4074_), .vdd(vdd), .B(raddr2_0_bF_buf70_), );
  OAI21X1 OAI21X1_1596 (.gnd(gnd), .A(_1138_), .Y(_4075_), .vdd(vdd), .B(raddr2_0_bF_buf69_), .C(_4074_), );
  NAND2X1 NAND2X1_706 (.gnd(gnd), .A(regs_24__0_), .Y(_4076_), .vdd(vdd), .B(raddr2_0_bF_buf68_), );
  OAI21X1 OAI21X1_1597 (.gnd(gnd), .A(_2417_), .Y(_4077_), .vdd(vdd), .B(raddr2_0_bF_buf67_), .C(_4076_), );
  MUX2X1 MUX2X1_306 (.gnd(gnd), .A(_4077_), .Y(_4078_), .vdd(vdd), .B(_4075_), .S(raddr2_1_bF_buf5_), );
  MUX2X1 MUX2X1_307 (.gnd(gnd), .A(_4078_), .Y(_4079_), .vdd(vdd), .B(_4073_), .S(raddr2_2_bF_buf7_), );
  MUX2X1 MUX2X1_308 (.gnd(gnd), .A(_4079_), .Y(_4080_), .vdd(vdd), .B(_4070_), .S(_4033__bF_buf6), );
  MUX2X1 MUX2X1_309 (.gnd(gnd), .A(_4058_), .Y(_5512__0_), .vdd(vdd), .B(_4080_), .S(raddr2_4_bF_buf4_), );
  OAI21X1 OAI21X1_1598 (.gnd(gnd), .A(_2479_), .Y(_4081_), .vdd(vdd), .B(raddr2_0_bF_buf66_), .C(raddr2_1_bF_buf4_), );
  AOI21X1 AOI21X1_250 (.gnd(gnd), .A(regs_4__1_), .Y(_4082_), .vdd(vdd), .B(raddr2_0_bF_buf65_), .C(_4081_), );
  AND2X2 AND2X2_44 (.gnd(gnd), .A(regs_6__1_), .Y(_4083_), .vdd(vdd), .B(raddr2_0_bF_buf64_), );
  OAI21X1 OAI21X1_1599 (.gnd(gnd), .A(_2103_), .Y(_4084_), .vdd(vdd), .B(raddr2_0_bF_buf63_), .C(_4038__bF_buf5), );
  OAI21X1 OAI21X1_1600 (.gnd(gnd), .A(_4084_), .Y(_4085_), .vdd(vdd), .B(_4083_), .C(_4036__bF_buf5), );
  OAI21X1 OAI21X1_1601 (.gnd(gnd), .A(_2486_), .Y(_4086_), .vdd(vdd), .B(raddr2_0_bF_buf62_), .C(raddr2_1_bF_buf3_), );
  AOI21X1 AOI21X1_251 (.gnd(gnd), .A(regs_0__1_), .Y(_4087_), .vdd(vdd), .B(raddr2_0_bF_buf61_), .C(_4086_), );
  NOR2X1 NOR2X1_196 (.gnd(gnd), .A(raddr2_0_bF_buf60_), .Y(_4088_), .vdd(vdd), .B(_2483_), );
  NAND2X1 NAND2X1_707 (.gnd(gnd), .A(regs_2__1_), .Y(_4089_), .vdd(vdd), .B(raddr2_0_bF_buf59_), );
  NAND2X1 NAND2X1_708 (.gnd(gnd), .A(_4038__bF_buf4), .Y(_4090_), .vdd(vdd), .B(_4089_), );
  OAI21X1 OAI21X1_1602 (.gnd(gnd), .A(_4090_), .Y(_4091_), .vdd(vdd), .B(_4088_), .C(raddr2_2_bF_buf6_), );
  OAI22X1 OAI22X1_55 (.gnd(gnd), .A(_4087_), .Y(_4092_), .vdd(vdd), .B(_4091_), .C(_4085_), .D(_4082_), );
  NAND2X1 NAND2X1_709 (.gnd(gnd), .A(regs_10__1_), .Y(_4093_), .vdd(vdd), .B(raddr2_0_bF_buf58_), );
  OAI21X1 OAI21X1_1603 (.gnd(gnd), .A(_1904_), .Y(_4094_), .vdd(vdd), .B(raddr2_0_bF_buf57_), .C(_4093_), );
  NAND2X1 NAND2X1_710 (.gnd(gnd), .A(regs_8__1_), .Y(_4095_), .vdd(vdd), .B(raddr2_0_bF_buf56_), );
  OAI21X1 OAI21X1_1604 (.gnd(gnd), .A(_2002_), .Y(_4096_), .vdd(vdd), .B(raddr2_0_bF_buf55_), .C(_4095_), );
  MUX2X1 MUX2X1_310 (.gnd(gnd), .A(_4096_), .Y(_4097_), .vdd(vdd), .B(_4094_), .S(raddr2_1_bF_buf2_), );
  NAND2X1 NAND2X1_711 (.gnd(gnd), .A(regs_14__1_), .Y(_4098_), .vdd(vdd), .B(raddr2_0_bF_buf54_), );
  OAI21X1 OAI21X1_1605 (.gnd(gnd), .A(_1707_), .Y(_4099_), .vdd(vdd), .B(raddr2_0_bF_buf53_), .C(_4098_), );
  NAND2X1 NAND2X1_712 (.gnd(gnd), .A(regs_12__1_), .Y(_4100_), .vdd(vdd), .B(raddr2_0_bF_buf52_), );
  OAI21X1 OAI21X1_1606 (.gnd(gnd), .A(_1805_), .Y(_4101_), .vdd(vdd), .B(raddr2_0_bF_buf51_), .C(_4100_), );
  MUX2X1 MUX2X1_311 (.gnd(gnd), .A(_4101_), .Y(_4102_), .vdd(vdd), .B(_4099_), .S(raddr2_1_bF_buf1_), );
  MUX2X1 MUX2X1_312 (.gnd(gnd), .A(_4102_), .Y(_4103_), .vdd(vdd), .B(_4097_), .S(_4036__bF_buf4), );
  MUX2X1 MUX2X1_313 (.gnd(gnd), .A(_4103_), .Y(_4104_), .vdd(vdd), .B(_4092_), .S(_4033__bF_buf5), );
  OAI21X1 OAI21X1_1607 (.gnd(gnd), .A(_1607_), .Y(_4105_), .vdd(vdd), .B(raddr2_0_bF_buf50_), .C(raddr2_1_bF_buf0_), );
  AOI21X1 AOI21X1_252 (.gnd(gnd), .A(regs_16__1_), .Y(_4106_), .vdd(vdd), .B(raddr2_0_bF_buf49_), .C(_4105_), );
  NOR2X1 NOR2X1_197 (.gnd(gnd), .A(raddr2_0_bF_buf48_), .Y(_4107_), .vdd(vdd), .B(_1509_), );
  NAND2X1 NAND2X1_713 (.gnd(gnd), .A(regs_18__1_), .Y(_4108_), .vdd(vdd), .B(raddr2_0_bF_buf47_), );
  NAND2X1 NAND2X1_714 (.gnd(gnd), .A(_4038__bF_buf3), .Y(_4109_), .vdd(vdd), .B(_4108_), );
  OAI21X1 OAI21X1_1608 (.gnd(gnd), .A(_4109_), .Y(_4110_), .vdd(vdd), .B(_4107_), .C(raddr2_2_bF_buf5_), );
  OAI21X1 OAI21X1_1609 (.gnd(gnd), .A(_1410_), .Y(_4111_), .vdd(vdd), .B(raddr2_0_bF_buf46_), .C(raddr2_1_bF_buf14_bF_buf2_), );
  AOI21X1 AOI21X1_253 (.gnd(gnd), .A(regs_20__1_), .Y(_4112_), .vdd(vdd), .B(raddr2_0_bF_buf45_), .C(_4111_), );
  AND2X2 AND2X2_45 (.gnd(gnd), .A(regs_22__1_), .Y(_4113_), .vdd(vdd), .B(raddr2_0_bF_buf44_), );
  OAI21X1 OAI21X1_1610 (.gnd(gnd), .A(_1312_), .Y(_4114_), .vdd(vdd), .B(raddr2_0_bF_buf43_), .C(_4038__bF_buf2), );
  OAI21X1 OAI21X1_1611 (.gnd(gnd), .A(_4114_), .Y(_4115_), .vdd(vdd), .B(_4113_), .C(_4036__bF_buf3), );
  OAI22X1 OAI22X1_56 (.gnd(gnd), .A(_4106_), .Y(_4116_), .vdd(vdd), .B(_4110_), .C(_4115_), .D(_4112_), );
  NAND2X1 NAND2X1_715 (.gnd(gnd), .A(regs_28__1_), .Y(_4117_), .vdd(vdd), .B(raddr2_0_bF_buf42_), );
  OAI21X1 OAI21X1_1612 (.gnd(gnd), .A(_2465_), .Y(_4118_), .vdd(vdd), .B(raddr2_0_bF_buf41_), .C(_4117_), );
  MUX2X1 MUX2X1_314 (.gnd(gnd), .A(_4118_), .Y(_4119_), .vdd(vdd), .B(regs_30__1_), .S(raddr2_1_bF_buf13_bF_buf2_), );
  NAND2X1 NAND2X1_716 (.gnd(gnd), .A(regs_26__1_), .Y(_4120_), .vdd(vdd), .B(raddr2_0_bF_buf40_), );
  OAI21X1 OAI21X1_1613 (.gnd(gnd), .A(_1145_), .Y(_4121_), .vdd(vdd), .B(raddr2_0_bF_buf39_), .C(_4120_), );
  NAND2X1 NAND2X1_717 (.gnd(gnd), .A(regs_24__1_), .Y(_4122_), .vdd(vdd), .B(raddr2_0_bF_buf38_), );
  OAI21X1 OAI21X1_1614 (.gnd(gnd), .A(_2471_), .Y(_4123_), .vdd(vdd), .B(raddr2_0_bF_buf37_), .C(_4122_), );
  MUX2X1 MUX2X1_315 (.gnd(gnd), .A(_4123_), .Y(_4124_), .vdd(vdd), .B(_4121_), .S(raddr2_1_bF_buf12_bF_buf2_), );
  MUX2X1 MUX2X1_316 (.gnd(gnd), .A(_4124_), .Y(_4125_), .vdd(vdd), .B(_4119_), .S(raddr2_2_bF_buf4_), );
  MUX2X1 MUX2X1_317 (.gnd(gnd), .A(_4125_), .Y(_4126_), .vdd(vdd), .B(_4116_), .S(_4033__bF_buf4), );
  MUX2X1 MUX2X1_318 (.gnd(gnd), .A(_4104_), .Y(_5512__1_), .vdd(vdd), .B(_4126_), .S(raddr2_4_bF_buf3_), );
  NAND2X1 NAND2X1_718 (.gnd(gnd), .A(regs_22__2_), .Y(_4127_), .vdd(vdd), .B(raddr2_0_bF_buf36_), );
  OAI21X1 OAI21X1_1615 (.gnd(gnd), .A(_1314_), .Y(_4128_), .vdd(vdd), .B(raddr2_0_bF_buf35_), .C(_4127_), );
  NAND2X1 NAND2X1_719 (.gnd(gnd), .A(regs_20__2_), .Y(_4129_), .vdd(vdd), .B(raddr2_0_bF_buf34_), );
  OAI21X1 OAI21X1_1616 (.gnd(gnd), .A(_1412_), .Y(_4130_), .vdd(vdd), .B(raddr2_0_bF_buf33_), .C(_4129_), );
  MUX2X1 MUX2X1_319 (.gnd(gnd), .A(_4130_), .Y(_4131_), .vdd(vdd), .B(_4128_), .S(raddr2_1_bF_buf11_), );
  NAND2X1 NAND2X1_720 (.gnd(gnd), .A(_4036__bF_buf2), .Y(_4132_), .vdd(vdd), .B(_4131_), );
  NAND2X1 NAND2X1_721 (.gnd(gnd), .A(regs_18__2_), .Y(_4133_), .vdd(vdd), .B(raddr2_0_bF_buf32_), );
  OAI21X1 OAI21X1_1617 (.gnd(gnd), .A(_1511_), .Y(_4134_), .vdd(vdd), .B(raddr2_0_bF_buf31_), .C(_4133_), );
  NAND2X1 NAND2X1_722 (.gnd(gnd), .A(regs_16__2_), .Y(_4135_), .vdd(vdd), .B(raddr2_0_bF_buf30_), );
  OAI21X1 OAI21X1_1618 (.gnd(gnd), .A(_1609_), .Y(_4136_), .vdd(vdd), .B(raddr2_0_bF_buf29_), .C(_4135_), );
  MUX2X1 MUX2X1_320 (.gnd(gnd), .A(_4136_), .Y(_4137_), .vdd(vdd), .B(_4134_), .S(raddr2_1_bF_buf10_), );
  AOI21X1 AOI21X1_254 (.gnd(gnd), .A(raddr2_2_bF_buf3_), .Y(_4138_), .vdd(vdd), .B(_4137_), .C(_4033__bF_buf3), );
  OAI21X1 OAI21X1_1619 (.gnd(gnd), .A(_1147_), .Y(_4139_), .vdd(vdd), .B(raddr2_0_bF_buf28_), .C(raddr2_2_bF_buf2_), );
  AOI21X1 AOI21X1_255 (.gnd(gnd), .A(regs_26__2_), .Y(_4140_), .vdd(vdd), .B(raddr2_0_bF_buf27_), .C(_4139_), );
  OAI21X1 OAI21X1_1620 (.gnd(gnd), .A(regs_30__2_), .Y(_4141_), .vdd(vdd), .B(raddr2_2_bF_buf1_), .C(_4038__bF_buf1), );
  OAI21X1 OAI21X1_1621 (.gnd(gnd), .A(_2518_), .Y(_4142_), .vdd(vdd), .B(raddr2_0_bF_buf26_), .C(raddr2_2_bF_buf0_), );
  AOI21X1 AOI21X1_256 (.gnd(gnd), .A(regs_24__2_), .Y(_4143_), .vdd(vdd), .B(raddr2_0_bF_buf25_), .C(_4142_), );
  NOR2X1 NOR2X1_198 (.gnd(gnd), .A(raddr2_0_bF_buf24_), .Y(_4144_), .vdd(vdd), .B(_2521_), );
  NAND2X1 NAND2X1_723 (.gnd(gnd), .A(regs_28__2_), .Y(_4145_), .vdd(vdd), .B(raddr2_0_bF_buf23_), );
  NAND2X1 NAND2X1_724 (.gnd(gnd), .A(_4036__bF_buf1), .Y(_4146_), .vdd(vdd), .B(_4145_), );
  OAI21X1 OAI21X1_1622 (.gnd(gnd), .A(_4146_), .Y(_4147_), .vdd(vdd), .B(_4144_), .C(raddr2_1_bF_buf9_), );
  OAI22X1 OAI22X1_57 (.gnd(gnd), .A(_4140_), .Y(_4148_), .vdd(vdd), .B(_4141_), .C(_4147_), .D(_4143_), );
  AOI22X1 AOI22X1_13 (.gnd(gnd), .A(_4148_), .Y(_4149_), .vdd(vdd), .B(_4033__bF_buf2), .C(_4132_), .D(_4138_), );
  OAI21X1 OAI21X1_1623 (.gnd(gnd), .A(_2530_), .Y(_4150_), .vdd(vdd), .B(raddr2_0_bF_buf22_), .C(raddr2_1_bF_buf8_), );
  AOI21X1 AOI21X1_257 (.gnd(gnd), .A(regs_4__2_), .Y(_4151_), .vdd(vdd), .B(raddr2_0_bF_buf21_), .C(_4150_), );
  AND2X2 AND2X2_46 (.gnd(gnd), .A(regs_6__2_), .Y(_4152_), .vdd(vdd), .B(raddr2_0_bF_buf20_), );
  OAI21X1 OAI21X1_1624 (.gnd(gnd), .A(_2105_), .Y(_4153_), .vdd(vdd), .B(raddr2_0_bF_buf19_), .C(_4038__bF_buf0), );
  OAI21X1 OAI21X1_1625 (.gnd(gnd), .A(_4153_), .Y(_4154_), .vdd(vdd), .B(_4152_), .C(_4036__bF_buf0), );
  OAI21X1 OAI21X1_1626 (.gnd(gnd), .A(_2537_), .Y(_4155_), .vdd(vdd), .B(raddr2_0_bF_buf18_), .C(raddr2_1_bF_buf7_), );
  AOI21X1 AOI21X1_258 (.gnd(gnd), .A(regs_0__2_), .Y(_4156_), .vdd(vdd), .B(raddr2_0_bF_buf17_), .C(_4155_), );
  NOR2X1 NOR2X1_199 (.gnd(gnd), .A(raddr2_0_bF_buf16_), .Y(_4157_), .vdd(vdd), .B(_2534_), );
  NAND2X1 NAND2X1_725 (.gnd(gnd), .A(regs_2__2_), .Y(_4158_), .vdd(vdd), .B(raddr2_0_bF_buf15_), );
  NAND2X1 NAND2X1_726 (.gnd(gnd), .A(_4038__bF_buf8), .Y(_4159_), .vdd(vdd), .B(_4158_), );
  OAI21X1 OAI21X1_1627 (.gnd(gnd), .A(_4159_), .Y(_4160_), .vdd(vdd), .B(_4157_), .C(raddr2_2_bF_buf10_), );
  OAI22X1 OAI22X1_58 (.gnd(gnd), .A(_4156_), .Y(_4161_), .vdd(vdd), .B(_4160_), .C(_4154_), .D(_4151_), );
  NAND2X1 NAND2X1_727 (.gnd(gnd), .A(regs_10__2_), .Y(_4162_), .vdd(vdd), .B(raddr2_0_bF_buf14_), );
  OAI21X1 OAI21X1_1628 (.gnd(gnd), .A(_1906_), .Y(_4163_), .vdd(vdd), .B(raddr2_0_bF_buf13_), .C(_4162_), );
  NAND2X1 NAND2X1_728 (.gnd(gnd), .A(regs_8__2_), .Y(_4164_), .vdd(vdd), .B(raddr2_0_bF_buf12_), );
  OAI21X1 OAI21X1_1629 (.gnd(gnd), .A(_2004_), .Y(_4165_), .vdd(vdd), .B(raddr2_0_bF_buf11_), .C(_4164_), );
  MUX2X1 MUX2X1_321 (.gnd(gnd), .A(_4165_), .Y(_4166_), .vdd(vdd), .B(_4163_), .S(raddr2_1_bF_buf6_), );
  NAND2X1 NAND2X1_729 (.gnd(gnd), .A(regs_14__2_), .Y(_4167_), .vdd(vdd), .B(raddr2_0_bF_buf10_), );
  OAI21X1 OAI21X1_1630 (.gnd(gnd), .A(_1709_), .Y(_4168_), .vdd(vdd), .B(raddr2_0_bF_buf9_), .C(_4167_), );
  NAND2X1 NAND2X1_730 (.gnd(gnd), .A(regs_12__2_), .Y(_4169_), .vdd(vdd), .B(raddr2_0_bF_buf8_), );
  OAI21X1 OAI21X1_1631 (.gnd(gnd), .A(_1807_), .Y(_4170_), .vdd(vdd), .B(raddr2_0_bF_buf7_), .C(_4169_), );
  MUX2X1 MUX2X1_322 (.gnd(gnd), .A(_4170_), .Y(_4171_), .vdd(vdd), .B(_4168_), .S(raddr2_1_bF_buf5_), );
  MUX2X1 MUX2X1_323 (.gnd(gnd), .A(_4171_), .Y(_4172_), .vdd(vdd), .B(_4166_), .S(_4036__bF_buf8), );
  MUX2X1 MUX2X1_324 (.gnd(gnd), .A(_4172_), .Y(_4173_), .vdd(vdd), .B(_4161_), .S(_4033__bF_buf1), );
  MUX2X1 MUX2X1_325 (.gnd(gnd), .A(_4173_), .Y(_5512__2_), .vdd(vdd), .B(_4149_), .S(raddr2_4_bF_buf2_), );
  NAND2X1 NAND2X1_731 (.gnd(gnd), .A(regs_22__3_), .Y(_4174_), .vdd(vdd), .B(raddr2_0_bF_buf6_), );
  OAI21X1 OAI21X1_1632 (.gnd(gnd), .A(_1316_), .Y(_4175_), .vdd(vdd), .B(raddr2_0_bF_buf5_), .C(_4174_), );
  NAND2X1 NAND2X1_732 (.gnd(gnd), .A(regs_20__3_), .Y(_4176_), .vdd(vdd), .B(raddr2_0_bF_buf4_), );
  OAI21X1 OAI21X1_1633 (.gnd(gnd), .A(_1414_), .Y(_4177_), .vdd(vdd), .B(raddr2_0_bF_buf3_), .C(_4176_), );
  MUX2X1 MUX2X1_326 (.gnd(gnd), .A(_4177_), .Y(_4178_), .vdd(vdd), .B(_4175_), .S(raddr2_1_bF_buf4_), );
  NAND2X1 NAND2X1_733 (.gnd(gnd), .A(_4036__bF_buf7), .Y(_4179_), .vdd(vdd), .B(_4178_), );
  NAND2X1 NAND2X1_734 (.gnd(gnd), .A(regs_18__3_), .Y(_4180_), .vdd(vdd), .B(raddr2_0_bF_buf2_), );
  OAI21X1 OAI21X1_1634 (.gnd(gnd), .A(_1513_), .Y(_4181_), .vdd(vdd), .B(raddr2_0_bF_buf1_), .C(_4180_), );
  NAND2X1 NAND2X1_735 (.gnd(gnd), .A(regs_16__3_), .Y(_4182_), .vdd(vdd), .B(raddr2_0_bF_buf0_), );
  OAI21X1 OAI21X1_1635 (.gnd(gnd), .A(_1611_), .Y(_4183_), .vdd(vdd), .B(raddr2_0_bF_buf96_), .C(_4182_), );
  MUX2X1 MUX2X1_327 (.gnd(gnd), .A(_4183_), .Y(_4184_), .vdd(vdd), .B(_4181_), .S(raddr2_1_bF_buf3_), );
  AOI21X1 AOI21X1_259 (.gnd(gnd), .A(raddr2_2_bF_buf9_), .Y(_4185_), .vdd(vdd), .B(_4184_), .C(_4033__bF_buf0), );
  OAI21X1 OAI21X1_1636 (.gnd(gnd), .A(_1149_), .Y(_4186_), .vdd(vdd), .B(raddr2_0_bF_buf95_), .C(raddr2_2_bF_buf8_), );
  AOI21X1 AOI21X1_260 (.gnd(gnd), .A(regs_26__3_), .Y(_4187_), .vdd(vdd), .B(raddr2_0_bF_buf94_), .C(_4186_), );
  OAI21X1 OAI21X1_1637 (.gnd(gnd), .A(regs_30__3_), .Y(_4188_), .vdd(vdd), .B(raddr2_2_bF_buf7_), .C(_4038__bF_buf7), );
  OAI21X1 OAI21X1_1638 (.gnd(gnd), .A(_2599_), .Y(_4189_), .vdd(vdd), .B(raddr2_0_bF_buf93_), .C(raddr2_2_bF_buf6_), );
  AOI21X1 AOI21X1_261 (.gnd(gnd), .A(regs_24__3_), .Y(_4190_), .vdd(vdd), .B(raddr2_0_bF_buf92_), .C(_4189_), );
  NOR2X1 NOR2X1_200 (.gnd(gnd), .A(raddr2_0_bF_buf91_), .Y(_4191_), .vdd(vdd), .B(_2593_), );
  NAND2X1 NAND2X1_736 (.gnd(gnd), .A(regs_28__3_), .Y(_4192_), .vdd(vdd), .B(raddr2_0_bF_buf90_), );
  NAND2X1 NAND2X1_737 (.gnd(gnd), .A(_4036__bF_buf6), .Y(_4193_), .vdd(vdd), .B(_4192_), );
  OAI21X1 OAI21X1_1639 (.gnd(gnd), .A(_4193_), .Y(_4194_), .vdd(vdd), .B(_4191_), .C(raddr2_1_bF_buf2_), );
  OAI22X1 OAI22X1_59 (.gnd(gnd), .A(_4187_), .Y(_4195_), .vdd(vdd), .B(_4188_), .C(_4194_), .D(_4190_), );
  AOI22X1 AOI22X1_14 (.gnd(gnd), .A(_4195_), .Y(_4196_), .vdd(vdd), .B(_4033__bF_buf7), .C(_4179_), .D(_4185_), );
  OAI21X1 OAI21X1_1640 (.gnd(gnd), .A(_2554_), .Y(_4197_), .vdd(vdd), .B(raddr2_0_bF_buf89_), .C(raddr2_1_bF_buf1_), );
  AOI21X1 AOI21X1_262 (.gnd(gnd), .A(regs_4__3_), .Y(_4198_), .vdd(vdd), .B(raddr2_0_bF_buf88_), .C(_4197_), );
  AND2X2 AND2X2_47 (.gnd(gnd), .A(regs_6__3_), .Y(_4199_), .vdd(vdd), .B(raddr2_0_bF_buf87_), );
  OAI21X1 OAI21X1_1641 (.gnd(gnd), .A(_2107_), .Y(_4200_), .vdd(vdd), .B(raddr2_0_bF_buf86_), .C(_4038__bF_buf6), );
  OAI21X1 OAI21X1_1642 (.gnd(gnd), .A(_4200_), .Y(_4201_), .vdd(vdd), .B(_4199_), .C(_4036__bF_buf5), );
  OAI21X1 OAI21X1_1643 (.gnd(gnd), .A(_2560_), .Y(_4202_), .vdd(vdd), .B(raddr2_0_bF_buf85_), .C(raddr2_1_bF_buf0_), );
  AOI21X1 AOI21X1_263 (.gnd(gnd), .A(regs_0__3_), .Y(_4203_), .vdd(vdd), .B(raddr2_0_bF_buf84_), .C(_4202_), );
  NOR2X1 NOR2X1_201 (.gnd(gnd), .A(raddr2_0_bF_buf83_), .Y(_4204_), .vdd(vdd), .B(_2563_), );
  NAND2X1 NAND2X1_738 (.gnd(gnd), .A(regs_2__3_), .Y(_4205_), .vdd(vdd), .B(raddr2_0_bF_buf82_), );
  NAND2X1 NAND2X1_739 (.gnd(gnd), .A(_4038__bF_buf5), .Y(_4206_), .vdd(vdd), .B(_4205_), );
  OAI21X1 OAI21X1_1644 (.gnd(gnd), .A(_4206_), .Y(_4207_), .vdd(vdd), .B(_4204_), .C(raddr2_2_bF_buf5_), );
  OAI22X1 OAI22X1_60 (.gnd(gnd), .A(_4203_), .Y(_4208_), .vdd(vdd), .B(_4207_), .C(_4201_), .D(_4198_), );
  NAND2X1 NAND2X1_740 (.gnd(gnd), .A(regs_10__3_), .Y(_4209_), .vdd(vdd), .B(raddr2_0_bF_buf81_), );
  OAI21X1 OAI21X1_1645 (.gnd(gnd), .A(_1908_), .Y(_4210_), .vdd(vdd), .B(raddr2_0_bF_buf80_), .C(_4209_), );
  NAND2X1 NAND2X1_741 (.gnd(gnd), .A(regs_8__3_), .Y(_4211_), .vdd(vdd), .B(raddr2_0_bF_buf79_), );
  OAI21X1 OAI21X1_1646 (.gnd(gnd), .A(_2006_), .Y(_4212_), .vdd(vdd), .B(raddr2_0_bF_buf78_), .C(_4211_), );
  MUX2X1 MUX2X1_328 (.gnd(gnd), .A(_4212_), .Y(_4213_), .vdd(vdd), .B(_4210_), .S(raddr2_1_bF_buf14_bF_buf1_), );
  NAND2X1 NAND2X1_742 (.gnd(gnd), .A(regs_14__3_), .Y(_4214_), .vdd(vdd), .B(raddr2_0_bF_buf77_), );
  OAI21X1 OAI21X1_1647 (.gnd(gnd), .A(_1711_), .Y(_4215_), .vdd(vdd), .B(raddr2_0_bF_buf76_), .C(_4214_), );
  NAND2X1 NAND2X1_743 (.gnd(gnd), .A(regs_12__3_), .Y(_4216_), .vdd(vdd), .B(raddr2_0_bF_buf75_), );
  OAI21X1 OAI21X1_1648 (.gnd(gnd), .A(_1809_), .Y(_4217_), .vdd(vdd), .B(raddr2_0_bF_buf74_), .C(_4216_), );
  MUX2X1 MUX2X1_329 (.gnd(gnd), .A(_4217_), .Y(_4218_), .vdd(vdd), .B(_4215_), .S(raddr2_1_bF_buf13_bF_buf1_), );
  MUX2X1 MUX2X1_330 (.gnd(gnd), .A(_4218_), .Y(_4219_), .vdd(vdd), .B(_4213_), .S(_4036__bF_buf4), );
  MUX2X1 MUX2X1_331 (.gnd(gnd), .A(_4219_), .Y(_4220_), .vdd(vdd), .B(_4208_), .S(_4033__bF_buf6), );
  MUX2X1 MUX2X1_332 (.gnd(gnd), .A(_4220_), .Y(_5512__3_), .vdd(vdd), .B(_4196_), .S(raddr2_4_bF_buf1_), );
  OAI21X1 OAI21X1_1649 (.gnd(gnd), .A(_2605_), .Y(_4221_), .vdd(vdd), .B(raddr2_0_bF_buf73_), .C(raddr2_1_bF_buf12_bF_buf1_), );
  AOI21X1 AOI21X1_264 (.gnd(gnd), .A(regs_4__4_), .Y(_4222_), .vdd(vdd), .B(raddr2_0_bF_buf72_), .C(_4221_), );
  AND2X2 AND2X2_48 (.gnd(gnd), .A(regs_6__4_), .Y(_4223_), .vdd(vdd), .B(raddr2_0_bF_buf71_), );
  OAI21X1 OAI21X1_1650 (.gnd(gnd), .A(_2109_), .Y(_4224_), .vdd(vdd), .B(raddr2_0_bF_buf70_), .C(_4038__bF_buf4), );
  OAI21X1 OAI21X1_1651 (.gnd(gnd), .A(_4224_), .Y(_4225_), .vdd(vdd), .B(_4223_), .C(_4036__bF_buf3), );
  OAI21X1 OAI21X1_1652 (.gnd(gnd), .A(_2611_), .Y(_4226_), .vdd(vdd), .B(raddr2_0_bF_buf69_), .C(raddr2_1_bF_buf11_), );
  AOI21X1 AOI21X1_265 (.gnd(gnd), .A(regs_0__4_), .Y(_4227_), .vdd(vdd), .B(raddr2_0_bF_buf68_), .C(_4226_), );
  NOR2X1 NOR2X1_202 (.gnd(gnd), .A(raddr2_0_bF_buf67_), .Y(_4228_), .vdd(vdd), .B(_2614_), );
  NAND2X1 NAND2X1_744 (.gnd(gnd), .A(regs_2__4_), .Y(_4229_), .vdd(vdd), .B(raddr2_0_bF_buf66_), );
  NAND2X1 NAND2X1_745 (.gnd(gnd), .A(_4038__bF_buf3), .Y(_4230_), .vdd(vdd), .B(_4229_), );
  OAI21X1 OAI21X1_1653 (.gnd(gnd), .A(_4230_), .Y(_4231_), .vdd(vdd), .B(_4228_), .C(raddr2_2_bF_buf4_), );
  OAI22X1 OAI22X1_61 (.gnd(gnd), .A(_4227_), .Y(_4232_), .vdd(vdd), .B(_4231_), .C(_4225_), .D(_4222_), );
  NAND2X1 NAND2X1_746 (.gnd(gnd), .A(regs_10__4_), .Y(_4233_), .vdd(vdd), .B(raddr2_0_bF_buf65_), );
  OAI21X1 OAI21X1_1654 (.gnd(gnd), .A(_1910_), .Y(_4234_), .vdd(vdd), .B(raddr2_0_bF_buf64_), .C(_4233_), );
  NAND2X1 NAND2X1_747 (.gnd(gnd), .A(regs_8__4_), .Y(_4235_), .vdd(vdd), .B(raddr2_0_bF_buf63_), );
  OAI21X1 OAI21X1_1655 (.gnd(gnd), .A(_2008_), .Y(_4236_), .vdd(vdd), .B(raddr2_0_bF_buf62_), .C(_4235_), );
  MUX2X1 MUX2X1_333 (.gnd(gnd), .A(_4236_), .Y(_4237_), .vdd(vdd), .B(_4234_), .S(raddr2_1_bF_buf10_), );
  NAND2X1 NAND2X1_748 (.gnd(gnd), .A(regs_14__4_), .Y(_4238_), .vdd(vdd), .B(raddr2_0_bF_buf61_), );
  OAI21X1 OAI21X1_1656 (.gnd(gnd), .A(_1713_), .Y(_4239_), .vdd(vdd), .B(raddr2_0_bF_buf60_), .C(_4238_), );
  NAND2X1 NAND2X1_749 (.gnd(gnd), .A(regs_12__4_), .Y(_4240_), .vdd(vdd), .B(raddr2_0_bF_buf59_), );
  OAI21X1 OAI21X1_1657 (.gnd(gnd), .A(_1811_), .Y(_4241_), .vdd(vdd), .B(raddr2_0_bF_buf58_), .C(_4240_), );
  MUX2X1 MUX2X1_334 (.gnd(gnd), .A(_4241_), .Y(_4242_), .vdd(vdd), .B(_4239_), .S(raddr2_1_bF_buf9_), );
  MUX2X1 MUX2X1_335 (.gnd(gnd), .A(_4242_), .Y(_4243_), .vdd(vdd), .B(_4237_), .S(_4036__bF_buf2), );
  MUX2X1 MUX2X1_336 (.gnd(gnd), .A(_4243_), .Y(_4244_), .vdd(vdd), .B(_4232_), .S(_4033__bF_buf5), );
  OAI21X1 OAI21X1_1658 (.gnd(gnd), .A(_1613_), .Y(_4245_), .vdd(vdd), .B(raddr2_0_bF_buf57_), .C(raddr2_1_bF_buf8_), );
  AOI21X1 AOI21X1_266 (.gnd(gnd), .A(regs_16__4_), .Y(_4246_), .vdd(vdd), .B(raddr2_0_bF_buf56_), .C(_4245_), );
  NOR2X1 NOR2X1_203 (.gnd(gnd), .A(raddr2_0_bF_buf55_), .Y(_4247_), .vdd(vdd), .B(_1515_), );
  NAND2X1 NAND2X1_750 (.gnd(gnd), .A(regs_18__4_), .Y(_4248_), .vdd(vdd), .B(raddr2_0_bF_buf54_), );
  NAND2X1 NAND2X1_751 (.gnd(gnd), .A(_4038__bF_buf2), .Y(_4249_), .vdd(vdd), .B(_4248_), );
  OAI21X1 OAI21X1_1659 (.gnd(gnd), .A(_4249_), .Y(_4250_), .vdd(vdd), .B(_4247_), .C(raddr2_2_bF_buf3_), );
  OAI21X1 OAI21X1_1660 (.gnd(gnd), .A(_1416_), .Y(_4251_), .vdd(vdd), .B(raddr2_0_bF_buf53_), .C(raddr2_1_bF_buf7_), );
  AOI21X1 AOI21X1_267 (.gnd(gnd), .A(regs_20__4_), .Y(_4252_), .vdd(vdd), .B(raddr2_0_bF_buf52_), .C(_4251_), );
  AND2X2 AND2X2_49 (.gnd(gnd), .A(regs_22__4_), .Y(_4253_), .vdd(vdd), .B(raddr2_0_bF_buf51_), );
  OAI21X1 OAI21X1_1661 (.gnd(gnd), .A(_1318_), .Y(_4254_), .vdd(vdd), .B(raddr2_0_bF_buf50_), .C(_4038__bF_buf1), );
  OAI21X1 OAI21X1_1662 (.gnd(gnd), .A(_4254_), .Y(_4255_), .vdd(vdd), .B(_4253_), .C(_4036__bF_buf1), );
  OAI22X1 OAI22X1_62 (.gnd(gnd), .A(_4246_), .Y(_4256_), .vdd(vdd), .B(_4250_), .C(_4255_), .D(_4252_), );
  NAND2X1 NAND2X1_752 (.gnd(gnd), .A(regs_28__4_), .Y(_4257_), .vdd(vdd), .B(raddr2_0_bF_buf49_), );
  OAI21X1 OAI21X1_1663 (.gnd(gnd), .A(_2644_), .Y(_4258_), .vdd(vdd), .B(raddr2_0_bF_buf48_), .C(_4257_), );
  MUX2X1 MUX2X1_337 (.gnd(gnd), .A(_4258_), .Y(_4259_), .vdd(vdd), .B(regs_30__4_), .S(raddr2_1_bF_buf6_), );
  NAND2X1 NAND2X1_753 (.gnd(gnd), .A(regs_26__4_), .Y(_4260_), .vdd(vdd), .B(raddr2_0_bF_buf47_), );
  OAI21X1 OAI21X1_1664 (.gnd(gnd), .A(_1151_), .Y(_4261_), .vdd(vdd), .B(raddr2_0_bF_buf46_), .C(_4260_), );
  NAND2X1 NAND2X1_754 (.gnd(gnd), .A(regs_24__4_), .Y(_4262_), .vdd(vdd), .B(raddr2_0_bF_buf45_), );
  OAI21X1 OAI21X1_1665 (.gnd(gnd), .A(_2650_), .Y(_4263_), .vdd(vdd), .B(raddr2_0_bF_buf44_), .C(_4262_), );
  MUX2X1 MUX2X1_338 (.gnd(gnd), .A(_4263_), .Y(_4264_), .vdd(vdd), .B(_4261_), .S(raddr2_1_bF_buf5_), );
  MUX2X1 MUX2X1_339 (.gnd(gnd), .A(_4264_), .Y(_4265_), .vdd(vdd), .B(_4259_), .S(raddr2_2_bF_buf2_), );
  MUX2X1 MUX2X1_340 (.gnd(gnd), .A(_4265_), .Y(_4266_), .vdd(vdd), .B(_4256_), .S(_4033__bF_buf4), );
  MUX2X1 MUX2X1_341 (.gnd(gnd), .A(_4244_), .Y(_5512__4_), .vdd(vdd), .B(_4266_), .S(raddr2_4_bF_buf0_), );
  OAI21X1 OAI21X1_1666 (.gnd(gnd), .A(_1418_), .Y(_4267_), .vdd(vdd), .B(raddr2_0_bF_buf43_), .C(raddr2_1_bF_buf4_), );
  AOI21X1 AOI21X1_268 (.gnd(gnd), .A(regs_20__5_), .Y(_4268_), .vdd(vdd), .B(raddr2_0_bF_buf42_), .C(_4267_), );
  AND2X2 AND2X2_50 (.gnd(gnd), .A(regs_22__5_), .Y(_4269_), .vdd(vdd), .B(raddr2_0_bF_buf41_), );
  OAI21X1 OAI21X1_1667 (.gnd(gnd), .A(_1320_), .Y(_4270_), .vdd(vdd), .B(raddr2_0_bF_buf40_), .C(_4038__bF_buf0), );
  OAI21X1 OAI21X1_1668 (.gnd(gnd), .A(_4270_), .Y(_4271_), .vdd(vdd), .B(_4269_), .C(_4036__bF_buf0), );
  OAI21X1 OAI21X1_1669 (.gnd(gnd), .A(_1615_), .Y(_4272_), .vdd(vdd), .B(raddr2_0_bF_buf39_), .C(raddr2_1_bF_buf3_), );
  AOI21X1 AOI21X1_269 (.gnd(gnd), .A(regs_16__5_), .Y(_4273_), .vdd(vdd), .B(raddr2_0_bF_buf38_), .C(_4272_), );
  NOR2X1 NOR2X1_204 (.gnd(gnd), .A(raddr2_0_bF_buf37_), .Y(_4274_), .vdd(vdd), .B(_1517_), );
  NAND2X1 NAND2X1_755 (.gnd(gnd), .A(regs_18__5_), .Y(_4275_), .vdd(vdd), .B(raddr2_0_bF_buf36_), );
  NAND2X1 NAND2X1_756 (.gnd(gnd), .A(_4038__bF_buf8), .Y(_4276_), .vdd(vdd), .B(_4275_), );
  OAI21X1 OAI21X1_1670 (.gnd(gnd), .A(_4276_), .Y(_4277_), .vdd(vdd), .B(_4274_), .C(raddr2_2_bF_buf1_), );
  OAI22X1 OAI22X1_63 (.gnd(gnd), .A(_4273_), .Y(_4278_), .vdd(vdd), .B(_4277_), .C(_4271_), .D(_4268_), );
  NAND2X1 NAND2X1_757 (.gnd(gnd), .A(regs_28__5_), .Y(_4279_), .vdd(vdd), .B(raddr2_0_bF_buf35_), );
  OAI21X1 OAI21X1_1671 (.gnd(gnd), .A(_2668_), .Y(_4280_), .vdd(vdd), .B(raddr2_0_bF_buf34_), .C(_4279_), );
  MUX2X1 MUX2X1_342 (.gnd(gnd), .A(_4280_), .Y(_4281_), .vdd(vdd), .B(regs_30__5_), .S(raddr2_1_bF_buf2_), );
  NAND2X1 NAND2X1_758 (.gnd(gnd), .A(regs_26__5_), .Y(_4282_), .vdd(vdd), .B(raddr2_0_bF_buf33_), );
  OAI21X1 OAI21X1_1672 (.gnd(gnd), .A(_1153_), .Y(_4283_), .vdd(vdd), .B(raddr2_0_bF_buf32_), .C(_4282_), );
  NAND2X1 NAND2X1_759 (.gnd(gnd), .A(regs_24__5_), .Y(_4284_), .vdd(vdd), .B(raddr2_0_bF_buf31_), );
  OAI21X1 OAI21X1_1673 (.gnd(gnd), .A(_2674_), .Y(_4285_), .vdd(vdd), .B(raddr2_0_bF_buf30_), .C(_4284_), );
  MUX2X1 MUX2X1_343 (.gnd(gnd), .A(_4285_), .Y(_4286_), .vdd(vdd), .B(_4283_), .S(raddr2_1_bF_buf1_), );
  MUX2X1 MUX2X1_344 (.gnd(gnd), .A(_4286_), .Y(_4287_), .vdd(vdd), .B(_4281_), .S(raddr2_2_bF_buf0_), );
  MUX2X1 MUX2X1_345 (.gnd(gnd), .A(_4287_), .Y(_4288_), .vdd(vdd), .B(_4278_), .S(_4033__bF_buf3), );
  NAND2X1 NAND2X1_760 (.gnd(gnd), .A(regs_6__5_), .Y(_4289_), .vdd(vdd), .B(raddr2_0_bF_buf29_), );
  OAI21X1 OAI21X1_1674 (.gnd(gnd), .A(_2111_), .Y(_4290_), .vdd(vdd), .B(raddr2_0_bF_buf28_), .C(_4289_), );
  NAND2X1 NAND2X1_761 (.gnd(gnd), .A(regs_4__5_), .Y(_4291_), .vdd(vdd), .B(raddr2_0_bF_buf27_), );
  OAI21X1 OAI21X1_1675 (.gnd(gnd), .A(_2682_), .Y(_4292_), .vdd(vdd), .B(raddr2_0_bF_buf26_), .C(_4291_), );
  MUX2X1 MUX2X1_346 (.gnd(gnd), .A(_4292_), .Y(_4293_), .vdd(vdd), .B(_4290_), .S(raddr2_1_bF_buf0_), );
  NAND2X1 NAND2X1_762 (.gnd(gnd), .A(regs_2__5_), .Y(_4294_), .vdd(vdd), .B(raddr2_0_bF_buf25_), );
  OAI21X1 OAI21X1_1676 (.gnd(gnd), .A(_2686_), .Y(_4295_), .vdd(vdd), .B(raddr2_0_bF_buf24_), .C(_4294_), );
  NAND2X1 NAND2X1_763 (.gnd(gnd), .A(regs_0__5_), .Y(_4296_), .vdd(vdd), .B(raddr2_0_bF_buf23_), );
  OAI21X1 OAI21X1_1677 (.gnd(gnd), .A(_2689_), .Y(_4297_), .vdd(vdd), .B(raddr2_0_bF_buf22_), .C(_4296_), );
  MUX2X1 MUX2X1_347 (.gnd(gnd), .A(_4297_), .Y(_4298_), .vdd(vdd), .B(_4295_), .S(raddr2_1_bF_buf14_bF_buf0_), );
  MUX2X1 MUX2X1_348 (.gnd(gnd), .A(_4298_), .Y(_4299_), .vdd(vdd), .B(_4293_), .S(raddr2_2_bF_buf10_), );
  NAND2X1 NAND2X1_764 (.gnd(gnd), .A(regs_14__5_), .Y(_4300_), .vdd(vdd), .B(raddr2_0_bF_buf21_), );
  OAI21X1 OAI21X1_1678 (.gnd(gnd), .A(_1715_), .Y(_4301_), .vdd(vdd), .B(raddr2_0_bF_buf20_), .C(_4300_), );
  NAND2X1 NAND2X1_765 (.gnd(gnd), .A(regs_12__5_), .Y(_4302_), .vdd(vdd), .B(raddr2_0_bF_buf19_), );
  OAI21X1 OAI21X1_1679 (.gnd(gnd), .A(_1813_), .Y(_4303_), .vdd(vdd), .B(raddr2_0_bF_buf18_), .C(_4302_), );
  MUX2X1 MUX2X1_349 (.gnd(gnd), .A(_4303_), .Y(_4304_), .vdd(vdd), .B(_4301_), .S(raddr2_1_bF_buf13_bF_buf0_), );
  NAND2X1 NAND2X1_766 (.gnd(gnd), .A(regs_10__5_), .Y(_4305_), .vdd(vdd), .B(raddr2_0_bF_buf17_), );
  OAI21X1 OAI21X1_1680 (.gnd(gnd), .A(_1912_), .Y(_4306_), .vdd(vdd), .B(raddr2_0_bF_buf16_), .C(_4305_), );
  NAND2X1 NAND2X1_767 (.gnd(gnd), .A(regs_8__5_), .Y(_4307_), .vdd(vdd), .B(raddr2_0_bF_buf15_), );
  OAI21X1 OAI21X1_1681 (.gnd(gnd), .A(_2010_), .Y(_4308_), .vdd(vdd), .B(raddr2_0_bF_buf14_), .C(_4307_), );
  MUX2X1 MUX2X1_350 (.gnd(gnd), .A(_4308_), .Y(_4309_), .vdd(vdd), .B(_4306_), .S(raddr2_1_bF_buf12_bF_buf0_), );
  MUX2X1 MUX2X1_351 (.gnd(gnd), .A(_4309_), .Y(_4310_), .vdd(vdd), .B(_4304_), .S(raddr2_2_bF_buf9_), );
  MUX2X1 MUX2X1_352 (.gnd(gnd), .A(_4310_), .Y(_4311_), .vdd(vdd), .B(_4299_), .S(_4033__bF_buf2), );
  MUX2X1 MUX2X1_353 (.gnd(gnd), .A(_4311_), .Y(_5512__5_), .vdd(vdd), .B(_4288_), .S(raddr2_4_bF_buf4_), );
  OAI21X1 OAI21X1_1682 (.gnd(gnd), .A(_1420_), .Y(_4312_), .vdd(vdd), .B(raddr2_0_bF_buf13_), .C(raddr2_1_bF_buf11_), );
  AOI21X1 AOI21X1_270 (.gnd(gnd), .A(regs_20__6_), .Y(_4313_), .vdd(vdd), .B(raddr2_0_bF_buf12_), .C(_4312_), );
  AND2X2 AND2X2_51 (.gnd(gnd), .A(regs_22__6_), .Y(_4314_), .vdd(vdd), .B(raddr2_0_bF_buf11_), );
  OAI21X1 OAI21X1_1683 (.gnd(gnd), .A(_1322_), .Y(_4315_), .vdd(vdd), .B(raddr2_0_bF_buf10_), .C(_4038__bF_buf7), );
  OAI21X1 OAI21X1_1684 (.gnd(gnd), .A(_4315_), .Y(_4316_), .vdd(vdd), .B(_4314_), .C(_4036__bF_buf8), );
  OAI21X1 OAI21X1_1685 (.gnd(gnd), .A(_1617_), .Y(_4317_), .vdd(vdd), .B(raddr2_0_bF_buf9_), .C(raddr2_1_bF_buf10_), );
  AOI21X1 AOI21X1_271 (.gnd(gnd), .A(regs_16__6_), .Y(_4318_), .vdd(vdd), .B(raddr2_0_bF_buf8_), .C(_4317_), );
  NOR2X1 NOR2X1_205 (.gnd(gnd), .A(raddr2_0_bF_buf7_), .Y(_4319_), .vdd(vdd), .B(_1519_), );
  NAND2X1 NAND2X1_768 (.gnd(gnd), .A(regs_18__6_), .Y(_4320_), .vdd(vdd), .B(raddr2_0_bF_buf6_), );
  NAND2X1 NAND2X1_769 (.gnd(gnd), .A(_4038__bF_buf6), .Y(_4321_), .vdd(vdd), .B(_4320_), );
  OAI21X1 OAI21X1_1686 (.gnd(gnd), .A(_4321_), .Y(_4322_), .vdd(vdd), .B(_4319_), .C(raddr2_2_bF_buf8_), );
  OAI22X1 OAI22X1_64 (.gnd(gnd), .A(_4318_), .Y(_4323_), .vdd(vdd), .B(_4322_), .C(_4316_), .D(_4313_), );
  NAND2X1 NAND2X1_770 (.gnd(gnd), .A(regs_28__6_), .Y(_4324_), .vdd(vdd), .B(raddr2_0_bF_buf5_), );
  OAI21X1 OAI21X1_1687 (.gnd(gnd), .A(_2718_), .Y(_4325_), .vdd(vdd), .B(raddr2_0_bF_buf4_), .C(_4324_), );
  MUX2X1 MUX2X1_354 (.gnd(gnd), .A(_4325_), .Y(_4326_), .vdd(vdd), .B(regs_30__6_), .S(raddr2_1_bF_buf9_), );
  NAND2X1 NAND2X1_771 (.gnd(gnd), .A(regs_26__6_), .Y(_4327_), .vdd(vdd), .B(raddr2_0_bF_buf3_), );
  OAI21X1 OAI21X1_1688 (.gnd(gnd), .A(_1155_), .Y(_4328_), .vdd(vdd), .B(raddr2_0_bF_buf2_), .C(_4327_), );
  NAND2X1 NAND2X1_772 (.gnd(gnd), .A(regs_24__6_), .Y(_4329_), .vdd(vdd), .B(raddr2_0_bF_buf1_), );
  OAI21X1 OAI21X1_1689 (.gnd(gnd), .A(_2724_), .Y(_4330_), .vdd(vdd), .B(raddr2_0_bF_buf0_), .C(_4329_), );
  MUX2X1 MUX2X1_355 (.gnd(gnd), .A(_4330_), .Y(_4331_), .vdd(vdd), .B(_4328_), .S(raddr2_1_bF_buf8_), );
  MUX2X1 MUX2X1_356 (.gnd(gnd), .A(_4331_), .Y(_4332_), .vdd(vdd), .B(_4326_), .S(raddr2_2_bF_buf7_), );
  MUX2X1 MUX2X1_357 (.gnd(gnd), .A(_4332_), .Y(_4333_), .vdd(vdd), .B(_4323_), .S(_4033__bF_buf1), );
  NAND2X1 NAND2X1_773 (.gnd(gnd), .A(regs_6__6_), .Y(_4334_), .vdd(vdd), .B(raddr2_0_bF_buf96_), );
  OAI21X1 OAI21X1_1690 (.gnd(gnd), .A(_2113_), .Y(_4335_), .vdd(vdd), .B(raddr2_0_bF_buf95_), .C(_4334_), );
  NAND2X1 NAND2X1_774 (.gnd(gnd), .A(regs_4__6_), .Y(_4336_), .vdd(vdd), .B(raddr2_0_bF_buf94_), );
  OAI21X1 OAI21X1_1691 (.gnd(gnd), .A(_2732_), .Y(_4337_), .vdd(vdd), .B(raddr2_0_bF_buf93_), .C(_4336_), );
  MUX2X1 MUX2X1_358 (.gnd(gnd), .A(_4337_), .Y(_4338_), .vdd(vdd), .B(_4335_), .S(raddr2_1_bF_buf7_), );
  NAND2X1 NAND2X1_775 (.gnd(gnd), .A(regs_2__6_), .Y(_4339_), .vdd(vdd), .B(raddr2_0_bF_buf92_), );
  OAI21X1 OAI21X1_1692 (.gnd(gnd), .A(_2736_), .Y(_4340_), .vdd(vdd), .B(raddr2_0_bF_buf91_), .C(_4339_), );
  NAND2X1 NAND2X1_776 (.gnd(gnd), .A(regs_0__6_), .Y(_4341_), .vdd(vdd), .B(raddr2_0_bF_buf90_), );
  OAI21X1 OAI21X1_1693 (.gnd(gnd), .A(_2739_), .Y(_4342_), .vdd(vdd), .B(raddr2_0_bF_buf89_), .C(_4341_), );
  MUX2X1 MUX2X1_359 (.gnd(gnd), .A(_4342_), .Y(_4343_), .vdd(vdd), .B(_4340_), .S(raddr2_1_bF_buf6_), );
  MUX2X1 MUX2X1_360 (.gnd(gnd), .A(_4343_), .Y(_4344_), .vdd(vdd), .B(_4338_), .S(raddr2_2_bF_buf6_), );
  NAND2X1 NAND2X1_777 (.gnd(gnd), .A(regs_14__6_), .Y(_4345_), .vdd(vdd), .B(raddr2_0_bF_buf88_), );
  OAI21X1 OAI21X1_1694 (.gnd(gnd), .A(_1717_), .Y(_4346_), .vdd(vdd), .B(raddr2_0_bF_buf87_), .C(_4345_), );
  NAND2X1 NAND2X1_778 (.gnd(gnd), .A(regs_12__6_), .Y(_4347_), .vdd(vdd), .B(raddr2_0_bF_buf86_), );
  OAI21X1 OAI21X1_1695 (.gnd(gnd), .A(_1815_), .Y(_4348_), .vdd(vdd), .B(raddr2_0_bF_buf85_), .C(_4347_), );
  MUX2X1 MUX2X1_361 (.gnd(gnd), .A(_4348_), .Y(_4349_), .vdd(vdd), .B(_4346_), .S(raddr2_1_bF_buf5_), );
  NAND2X1 NAND2X1_779 (.gnd(gnd), .A(regs_10__6_), .Y(_4350_), .vdd(vdd), .B(raddr2_0_bF_buf84_), );
  OAI21X1 OAI21X1_1696 (.gnd(gnd), .A(_1914_), .Y(_4351_), .vdd(vdd), .B(raddr2_0_bF_buf83_), .C(_4350_), );
  NAND2X1 NAND2X1_780 (.gnd(gnd), .A(regs_8__6_), .Y(_4352_), .vdd(vdd), .B(raddr2_0_bF_buf82_), );
  OAI21X1 OAI21X1_1697 (.gnd(gnd), .A(_2012_), .Y(_4353_), .vdd(vdd), .B(raddr2_0_bF_buf81_), .C(_4352_), );
  MUX2X1 MUX2X1_362 (.gnd(gnd), .A(_4353_), .Y(_4354_), .vdd(vdd), .B(_4351_), .S(raddr2_1_bF_buf4_), );
  MUX2X1 MUX2X1_363 (.gnd(gnd), .A(_4354_), .Y(_4355_), .vdd(vdd), .B(_4349_), .S(raddr2_2_bF_buf5_), );
  MUX2X1 MUX2X1_364 (.gnd(gnd), .A(_4355_), .Y(_4356_), .vdd(vdd), .B(_4344_), .S(_4033__bF_buf0), );
  MUX2X1 MUX2X1_365 (.gnd(gnd), .A(_4356_), .Y(_5512__6_), .vdd(vdd), .B(_4333_), .S(raddr2_4_bF_buf3_), );
  NAND2X1 NAND2X1_781 (.gnd(gnd), .A(regs_22__7_), .Y(_4357_), .vdd(vdd), .B(raddr2_0_bF_buf80_), );
  OAI21X1 OAI21X1_1698 (.gnd(gnd), .A(_1324_), .Y(_4358_), .vdd(vdd), .B(raddr2_0_bF_buf79_), .C(_4357_), );
  NAND2X1 NAND2X1_782 (.gnd(gnd), .A(regs_20__7_), .Y(_4359_), .vdd(vdd), .B(raddr2_0_bF_buf78_), );
  OAI21X1 OAI21X1_1699 (.gnd(gnd), .A(_1422_), .Y(_4360_), .vdd(vdd), .B(raddr2_0_bF_buf77_), .C(_4359_), );
  MUX2X1 MUX2X1_366 (.gnd(gnd), .A(_4360_), .Y(_4361_), .vdd(vdd), .B(_4358_), .S(raddr2_1_bF_buf3_), );
  NAND2X1 NAND2X1_783 (.gnd(gnd), .A(_4036__bF_buf7), .Y(_4362_), .vdd(vdd), .B(_4361_), );
  NAND2X1 NAND2X1_784 (.gnd(gnd), .A(regs_18__7_), .Y(_4363_), .vdd(vdd), .B(raddr2_0_bF_buf76_), );
  OAI21X1 OAI21X1_1700 (.gnd(gnd), .A(_1521_), .Y(_4364_), .vdd(vdd), .B(raddr2_0_bF_buf75_), .C(_4363_), );
  NAND2X1 NAND2X1_785 (.gnd(gnd), .A(regs_16__7_), .Y(_4365_), .vdd(vdd), .B(raddr2_0_bF_buf74_), );
  OAI21X1 OAI21X1_1701 (.gnd(gnd), .A(_1619_), .Y(_4366_), .vdd(vdd), .B(raddr2_0_bF_buf73_), .C(_4365_), );
  MUX2X1 MUX2X1_367 (.gnd(gnd), .A(_4366_), .Y(_4367_), .vdd(vdd), .B(_4364_), .S(raddr2_1_bF_buf2_), );
  AOI21X1 AOI21X1_272 (.gnd(gnd), .A(raddr2_2_bF_buf4_), .Y(_4368_), .vdd(vdd), .B(_4367_), .C(_4033__bF_buf7), );
  OAI21X1 OAI21X1_1702 (.gnd(gnd), .A(_1157_), .Y(_4369_), .vdd(vdd), .B(raddr2_0_bF_buf72_), .C(raddr2_2_bF_buf3_), );
  AOI21X1 AOI21X1_273 (.gnd(gnd), .A(regs_26__7_), .Y(_4370_), .vdd(vdd), .B(raddr2_0_bF_buf71_), .C(_4369_), );
  OAI21X1 OAI21X1_1703 (.gnd(gnd), .A(regs_30__7_), .Y(_4371_), .vdd(vdd), .B(raddr2_2_bF_buf2_), .C(_4038__bF_buf5), );
  OAI21X1 OAI21X1_1704 (.gnd(gnd), .A(_2771_), .Y(_4372_), .vdd(vdd), .B(raddr2_0_bF_buf70_), .C(raddr2_2_bF_buf1_), );
  AOI21X1 AOI21X1_274 (.gnd(gnd), .A(regs_24__7_), .Y(_4373_), .vdd(vdd), .B(raddr2_0_bF_buf69_), .C(_4372_), );
  NOR2X1 NOR2X1_206 (.gnd(gnd), .A(raddr2_0_bF_buf68_), .Y(_4374_), .vdd(vdd), .B(_2774_), );
  NAND2X1 NAND2X1_786 (.gnd(gnd), .A(regs_28__7_), .Y(_4375_), .vdd(vdd), .B(raddr2_0_bF_buf67_), );
  NAND2X1 NAND2X1_787 (.gnd(gnd), .A(_4036__bF_buf6), .Y(_4376_), .vdd(vdd), .B(_4375_), );
  OAI21X1 OAI21X1_1705 (.gnd(gnd), .A(_4376_), .Y(_4377_), .vdd(vdd), .B(_4374_), .C(raddr2_1_bF_buf1_), );
  OAI22X1 OAI22X1_65 (.gnd(gnd), .A(_4370_), .Y(_4378_), .vdd(vdd), .B(_4371_), .C(_4377_), .D(_4373_), );
  AOI22X1 AOI22X1_15 (.gnd(gnd), .A(_4378_), .Y(_4379_), .vdd(vdd), .B(_4033__bF_buf6), .C(_4362_), .D(_4368_), );
  OAI21X1 OAI21X1_1706 (.gnd(gnd), .A(_2781_), .Y(_4380_), .vdd(vdd), .B(raddr2_0_bF_buf66_), .C(raddr2_1_bF_buf0_), );
  AOI21X1 AOI21X1_275 (.gnd(gnd), .A(regs_4__7_), .Y(_4381_), .vdd(vdd), .B(raddr2_0_bF_buf65_), .C(_4380_), );
  AND2X2 AND2X2_52 (.gnd(gnd), .A(regs_6__7_), .Y(_4382_), .vdd(vdd), .B(raddr2_0_bF_buf64_), );
  OAI21X1 OAI21X1_1707 (.gnd(gnd), .A(_2115_), .Y(_4383_), .vdd(vdd), .B(raddr2_0_bF_buf63_), .C(_4038__bF_buf4), );
  OAI21X1 OAI21X1_1708 (.gnd(gnd), .A(_4383_), .Y(_4384_), .vdd(vdd), .B(_4382_), .C(_4036__bF_buf5), );
  OAI21X1 OAI21X1_1709 (.gnd(gnd), .A(_2787_), .Y(_4385_), .vdd(vdd), .B(raddr2_0_bF_buf62_), .C(raddr2_1_bF_buf14_bF_buf3_), );
  AOI21X1 AOI21X1_276 (.gnd(gnd), .A(regs_0__7_), .Y(_4386_), .vdd(vdd), .B(raddr2_0_bF_buf61_), .C(_4385_), );
  NOR2X1 NOR2X1_207 (.gnd(gnd), .A(raddr2_0_bF_buf60_), .Y(_4387_), .vdd(vdd), .B(_2790_), );
  NAND2X1 NAND2X1_788 (.gnd(gnd), .A(regs_2__7_), .Y(_4388_), .vdd(vdd), .B(raddr2_0_bF_buf59_), );
  NAND2X1 NAND2X1_789 (.gnd(gnd), .A(_4038__bF_buf3), .Y(_4389_), .vdd(vdd), .B(_4388_), );
  OAI21X1 OAI21X1_1710 (.gnd(gnd), .A(_4389_), .Y(_4390_), .vdd(vdd), .B(_4387_), .C(raddr2_2_bF_buf0_), );
  OAI22X1 OAI22X1_66 (.gnd(gnd), .A(_4386_), .Y(_4391_), .vdd(vdd), .B(_4390_), .C(_4384_), .D(_4381_), );
  NAND2X1 NAND2X1_790 (.gnd(gnd), .A(regs_10__7_), .Y(_4392_), .vdd(vdd), .B(raddr2_0_bF_buf58_), );
  OAI21X1 OAI21X1_1711 (.gnd(gnd), .A(_1916_), .Y(_4393_), .vdd(vdd), .B(raddr2_0_bF_buf57_), .C(_4392_), );
  NAND2X1 NAND2X1_791 (.gnd(gnd), .A(regs_8__7_), .Y(_4394_), .vdd(vdd), .B(raddr2_0_bF_buf56_), );
  OAI21X1 OAI21X1_1712 (.gnd(gnd), .A(_2014_), .Y(_4395_), .vdd(vdd), .B(raddr2_0_bF_buf55_), .C(_4394_), );
  MUX2X1 MUX2X1_368 (.gnd(gnd), .A(_4395_), .Y(_4396_), .vdd(vdd), .B(_4393_), .S(raddr2_1_bF_buf13_bF_buf3_), );
  NAND2X1 NAND2X1_792 (.gnd(gnd), .A(regs_14__7_), .Y(_4397_), .vdd(vdd), .B(raddr2_0_bF_buf54_), );
  OAI21X1 OAI21X1_1713 (.gnd(gnd), .A(_1719_), .Y(_4398_), .vdd(vdd), .B(raddr2_0_bF_buf53_), .C(_4397_), );
  NAND2X1 NAND2X1_793 (.gnd(gnd), .A(regs_12__7_), .Y(_4399_), .vdd(vdd), .B(raddr2_0_bF_buf52_), );
  OAI21X1 OAI21X1_1714 (.gnd(gnd), .A(_1817_), .Y(_4400_), .vdd(vdd), .B(raddr2_0_bF_buf51_), .C(_4399_), );
  MUX2X1 MUX2X1_369 (.gnd(gnd), .A(_4400_), .Y(_4401_), .vdd(vdd), .B(_4398_), .S(raddr2_1_bF_buf12_bF_buf3_), );
  MUX2X1 MUX2X1_370 (.gnd(gnd), .A(_4401_), .Y(_4402_), .vdd(vdd), .B(_4396_), .S(_4036__bF_buf4), );
  MUX2X1 MUX2X1_371 (.gnd(gnd), .A(_4402_), .Y(_4403_), .vdd(vdd), .B(_4391_), .S(_4033__bF_buf5), );
  MUX2X1 MUX2X1_372 (.gnd(gnd), .A(_4403_), .Y(_5512__7_), .vdd(vdd), .B(_4379_), .S(raddr2_4_bF_buf2_), );
  OAI21X1 OAI21X1_1715 (.gnd(gnd), .A(_1424_), .Y(_4404_), .vdd(vdd), .B(raddr2_0_bF_buf50_), .C(raddr2_1_bF_buf11_), );
  AOI21X1 AOI21X1_277 (.gnd(gnd), .A(regs_20__8_), .Y(_4405_), .vdd(vdd), .B(raddr2_0_bF_buf49_), .C(_4404_), );
  AND2X2 AND2X2_53 (.gnd(gnd), .A(regs_22__8_), .Y(_4406_), .vdd(vdd), .B(raddr2_0_bF_buf48_), );
  OAI21X1 OAI21X1_1716 (.gnd(gnd), .A(_1326_), .Y(_4407_), .vdd(vdd), .B(raddr2_0_bF_buf47_), .C(_4038__bF_buf2), );
  OAI21X1 OAI21X1_1717 (.gnd(gnd), .A(_4407_), .Y(_4408_), .vdd(vdd), .B(_4406_), .C(_4036__bF_buf3), );
  OAI21X1 OAI21X1_1718 (.gnd(gnd), .A(_1621_), .Y(_4409_), .vdd(vdd), .B(raddr2_0_bF_buf46_), .C(raddr2_1_bF_buf10_), );
  AOI21X1 AOI21X1_278 (.gnd(gnd), .A(regs_16__8_), .Y(_4410_), .vdd(vdd), .B(raddr2_0_bF_buf45_), .C(_4409_), );
  NOR2X1 NOR2X1_208 (.gnd(gnd), .A(raddr2_0_bF_buf44_), .Y(_4411_), .vdd(vdd), .B(_1523_), );
  NAND2X1 NAND2X1_794 (.gnd(gnd), .A(regs_18__8_), .Y(_4412_), .vdd(vdd), .B(raddr2_0_bF_buf43_), );
  NAND2X1 NAND2X1_795 (.gnd(gnd), .A(_4038__bF_buf1), .Y(_4413_), .vdd(vdd), .B(_4412_), );
  OAI21X1 OAI21X1_1719 (.gnd(gnd), .A(_4413_), .Y(_4414_), .vdd(vdd), .B(_4411_), .C(raddr2_2_bF_buf10_), );
  OAI22X1 OAI22X1_67 (.gnd(gnd), .A(_4410_), .Y(_4415_), .vdd(vdd), .B(_4414_), .C(_4408_), .D(_4405_), );
  NAND2X1 NAND2X1_796 (.gnd(gnd), .A(regs_28__8_), .Y(_4416_), .vdd(vdd), .B(raddr2_0_bF_buf42_), );
  OAI21X1 OAI21X1_1720 (.gnd(gnd), .A(_2847_), .Y(_4417_), .vdd(vdd), .B(raddr2_0_bF_buf41_), .C(_4416_), );
  MUX2X1 MUX2X1_373 (.gnd(gnd), .A(_4417_), .Y(_4418_), .vdd(vdd), .B(regs_30__8_), .S(raddr2_1_bF_buf9_), );
  NAND2X1 NAND2X1_797 (.gnd(gnd), .A(regs_26__8_), .Y(_4419_), .vdd(vdd), .B(raddr2_0_bF_buf40_), );
  OAI21X1 OAI21X1_1721 (.gnd(gnd), .A(_1159_), .Y(_4420_), .vdd(vdd), .B(raddr2_0_bF_buf39_), .C(_4419_), );
  NAND2X1 NAND2X1_798 (.gnd(gnd), .A(regs_24__8_), .Y(_4421_), .vdd(vdd), .B(raddr2_0_bF_buf38_), );
  OAI21X1 OAI21X1_1722 (.gnd(gnd), .A(_2853_), .Y(_4422_), .vdd(vdd), .B(raddr2_0_bF_buf37_), .C(_4421_), );
  MUX2X1 MUX2X1_374 (.gnd(gnd), .A(_4422_), .Y(_4423_), .vdd(vdd), .B(_4420_), .S(raddr2_1_bF_buf8_), );
  MUX2X1 MUX2X1_375 (.gnd(gnd), .A(_4423_), .Y(_4424_), .vdd(vdd), .B(_4418_), .S(raddr2_2_bF_buf9_), );
  MUX2X1 MUX2X1_376 (.gnd(gnd), .A(_4424_), .Y(_4425_), .vdd(vdd), .B(_4415_), .S(_4033__bF_buf4), );
  NAND2X1 NAND2X1_799 (.gnd(gnd), .A(regs_6__8_), .Y(_4426_), .vdd(vdd), .B(raddr2_0_bF_buf36_), );
  OAI21X1 OAI21X1_1723 (.gnd(gnd), .A(_2117_), .Y(_4427_), .vdd(vdd), .B(raddr2_0_bF_buf35_), .C(_4426_), );
  NAND2X1 NAND2X1_800 (.gnd(gnd), .A(regs_4__8_), .Y(_4428_), .vdd(vdd), .B(raddr2_0_bF_buf34_), );
  OAI21X1 OAI21X1_1724 (.gnd(gnd), .A(_2808_), .Y(_4429_), .vdd(vdd), .B(raddr2_0_bF_buf33_), .C(_4428_), );
  MUX2X1 MUX2X1_377 (.gnd(gnd), .A(_4429_), .Y(_4430_), .vdd(vdd), .B(_4427_), .S(raddr2_1_bF_buf7_), );
  NAND2X1 NAND2X1_801 (.gnd(gnd), .A(regs_2__8_), .Y(_4431_), .vdd(vdd), .B(raddr2_0_bF_buf32_), );
  OAI21X1 OAI21X1_1725 (.gnd(gnd), .A(_2817_), .Y(_4432_), .vdd(vdd), .B(raddr2_0_bF_buf31_), .C(_4431_), );
  NAND2X1 NAND2X1_802 (.gnd(gnd), .A(regs_0__8_), .Y(_4433_), .vdd(vdd), .B(raddr2_0_bF_buf30_), );
  OAI21X1 OAI21X1_1726 (.gnd(gnd), .A(_2814_), .Y(_4434_), .vdd(vdd), .B(raddr2_0_bF_buf29_), .C(_4433_), );
  MUX2X1 MUX2X1_378 (.gnd(gnd), .A(_4434_), .Y(_4435_), .vdd(vdd), .B(_4432_), .S(raddr2_1_bF_buf6_), );
  MUX2X1 MUX2X1_379 (.gnd(gnd), .A(_4435_), .Y(_4436_), .vdd(vdd), .B(_4430_), .S(raddr2_2_bF_buf8_), );
  NAND2X1 NAND2X1_803 (.gnd(gnd), .A(regs_14__8_), .Y(_4437_), .vdd(vdd), .B(raddr2_0_bF_buf28_), );
  OAI21X1 OAI21X1_1727 (.gnd(gnd), .A(_1721_), .Y(_4438_), .vdd(vdd), .B(raddr2_0_bF_buf27_), .C(_4437_), );
  NAND2X1 NAND2X1_804 (.gnd(gnd), .A(regs_12__8_), .Y(_4439_), .vdd(vdd), .B(raddr2_0_bF_buf26_), );
  OAI21X1 OAI21X1_1728 (.gnd(gnd), .A(_1819_), .Y(_4440_), .vdd(vdd), .B(raddr2_0_bF_buf25_), .C(_4439_), );
  MUX2X1 MUX2X1_380 (.gnd(gnd), .A(_4440_), .Y(_4441_), .vdd(vdd), .B(_4438_), .S(raddr2_1_bF_buf5_), );
  NAND2X1 NAND2X1_805 (.gnd(gnd), .A(regs_10__8_), .Y(_4442_), .vdd(vdd), .B(raddr2_0_bF_buf24_), );
  OAI21X1 OAI21X1_1729 (.gnd(gnd), .A(_1918_), .Y(_4443_), .vdd(vdd), .B(raddr2_0_bF_buf23_), .C(_4442_), );
  NAND2X1 NAND2X1_806 (.gnd(gnd), .A(regs_8__8_), .Y(_4444_), .vdd(vdd), .B(raddr2_0_bF_buf22_), );
  OAI21X1 OAI21X1_1730 (.gnd(gnd), .A(_2016_), .Y(_4445_), .vdd(vdd), .B(raddr2_0_bF_buf21_), .C(_4444_), );
  MUX2X1 MUX2X1_381 (.gnd(gnd), .A(_4445_), .Y(_4446_), .vdd(vdd), .B(_4443_), .S(raddr2_1_bF_buf4_), );
  MUX2X1 MUX2X1_382 (.gnd(gnd), .A(_4446_), .Y(_4447_), .vdd(vdd), .B(_4441_), .S(raddr2_2_bF_buf7_), );
  MUX2X1 MUX2X1_383 (.gnd(gnd), .A(_4447_), .Y(_4448_), .vdd(vdd), .B(_4436_), .S(_4033__bF_buf3), );
  MUX2X1 MUX2X1_384 (.gnd(gnd), .A(_4448_), .Y(_5512__8_), .vdd(vdd), .B(_4425_), .S(raddr2_4_bF_buf1_), );
  NAND2X1 NAND2X1_807 (.gnd(gnd), .A(regs_22__9_), .Y(_4449_), .vdd(vdd), .B(raddr2_0_bF_buf20_), );
  OAI21X1 OAI21X1_1731 (.gnd(gnd), .A(_1328_), .Y(_4450_), .vdd(vdd), .B(raddr2_0_bF_buf19_), .C(_4449_), );
  NAND2X1 NAND2X1_808 (.gnd(gnd), .A(regs_20__9_), .Y(_4451_), .vdd(vdd), .B(raddr2_0_bF_buf18_), );
  OAI21X1 OAI21X1_1732 (.gnd(gnd), .A(_1426_), .Y(_4452_), .vdd(vdd), .B(raddr2_0_bF_buf17_), .C(_4451_), );
  MUX2X1 MUX2X1_385 (.gnd(gnd), .A(_4452_), .Y(_4453_), .vdd(vdd), .B(_4450_), .S(raddr2_1_bF_buf3_), );
  NAND2X1 NAND2X1_809 (.gnd(gnd), .A(_4036__bF_buf2), .Y(_4454_), .vdd(vdd), .B(_4453_), );
  NAND2X1 NAND2X1_810 (.gnd(gnd), .A(regs_18__9_), .Y(_4455_), .vdd(vdd), .B(raddr2_0_bF_buf16_), );
  OAI21X1 OAI21X1_1733 (.gnd(gnd), .A(_1525_), .Y(_4456_), .vdd(vdd), .B(raddr2_0_bF_buf15_), .C(_4455_), );
  NAND2X1 NAND2X1_811 (.gnd(gnd), .A(regs_16__9_), .Y(_4457_), .vdd(vdd), .B(raddr2_0_bF_buf14_), );
  OAI21X1 OAI21X1_1734 (.gnd(gnd), .A(_1623_), .Y(_4458_), .vdd(vdd), .B(raddr2_0_bF_buf13_), .C(_4457_), );
  MUX2X1 MUX2X1_386 (.gnd(gnd), .A(_4458_), .Y(_4459_), .vdd(vdd), .B(_4456_), .S(raddr2_1_bF_buf2_), );
  AOI21X1 AOI21X1_279 (.gnd(gnd), .A(raddr2_2_bF_buf6_), .Y(_4460_), .vdd(vdd), .B(_4459_), .C(_4033__bF_buf2), );
  OAI21X1 OAI21X1_1735 (.gnd(gnd), .A(_1161_), .Y(_4461_), .vdd(vdd), .B(raddr2_0_bF_buf12_), .C(raddr2_2_bF_buf5_), );
  AOI21X1 AOI21X1_280 (.gnd(gnd), .A(regs_26__9_), .Y(_4462_), .vdd(vdd), .B(raddr2_0_bF_buf11_), .C(_4461_), );
  OAI21X1 OAI21X1_1736 (.gnd(gnd), .A(regs_30__9_), .Y(_4463_), .vdd(vdd), .B(raddr2_2_bF_buf4_), .C(_4038__bF_buf0), );
  OAI21X1 OAI21X1_1737 (.gnd(gnd), .A(_2874_), .Y(_4464_), .vdd(vdd), .B(raddr2_0_bF_buf10_), .C(raddr2_2_bF_buf3_), );
  AOI21X1 AOI21X1_281 (.gnd(gnd), .A(regs_24__9_), .Y(_4465_), .vdd(vdd), .B(raddr2_0_bF_buf9_), .C(_4464_), );
  NOR2X1 NOR2X1_209 (.gnd(gnd), .A(raddr2_0_bF_buf8_), .Y(_4466_), .vdd(vdd), .B(_2877_), );
  NAND2X1 NAND2X1_812 (.gnd(gnd), .A(regs_28__9_), .Y(_4467_), .vdd(vdd), .B(raddr2_0_bF_buf7_), );
  NAND2X1 NAND2X1_813 (.gnd(gnd), .A(_4036__bF_buf1), .Y(_4468_), .vdd(vdd), .B(_4467_), );
  OAI21X1 OAI21X1_1738 (.gnd(gnd), .A(_4468_), .Y(_4469_), .vdd(vdd), .B(_4466_), .C(raddr2_1_bF_buf1_), );
  OAI22X1 OAI22X1_68 (.gnd(gnd), .A(_4462_), .Y(_4470_), .vdd(vdd), .B(_4463_), .C(_4469_), .D(_4465_), );
  AOI22X1 AOI22X1_16 (.gnd(gnd), .A(_4470_), .Y(_4471_), .vdd(vdd), .B(_4033__bF_buf1), .C(_4454_), .D(_4460_), );
  OAI21X1 OAI21X1_1739 (.gnd(gnd), .A(_2886_), .Y(_4472_), .vdd(vdd), .B(raddr2_0_bF_buf6_), .C(raddr2_1_bF_buf0_), );
  AOI21X1 AOI21X1_282 (.gnd(gnd), .A(regs_4__9_), .Y(_4473_), .vdd(vdd), .B(raddr2_0_bF_buf5_), .C(_4472_), );
  AND2X2 AND2X2_54 (.gnd(gnd), .A(regs_6__9_), .Y(_4474_), .vdd(vdd), .B(raddr2_0_bF_buf4_), );
  OAI21X1 OAI21X1_1740 (.gnd(gnd), .A(_2119_), .Y(_4475_), .vdd(vdd), .B(raddr2_0_bF_buf3_), .C(_4038__bF_buf8), );
  OAI21X1 OAI21X1_1741 (.gnd(gnd), .A(_4475_), .Y(_4476_), .vdd(vdd), .B(_4474_), .C(_4036__bF_buf0), );
  OAI21X1 OAI21X1_1742 (.gnd(gnd), .A(_2893_), .Y(_4477_), .vdd(vdd), .B(raddr2_0_bF_buf2_), .C(raddr2_1_bF_buf14_bF_buf2_), );
  AOI21X1 AOI21X1_283 (.gnd(gnd), .A(regs_0__9_), .Y(_4478_), .vdd(vdd), .B(raddr2_0_bF_buf1_), .C(_4477_), );
  NOR2X1 NOR2X1_210 (.gnd(gnd), .A(raddr2_0_bF_buf0_), .Y(_4479_), .vdd(vdd), .B(_2890_), );
  NAND2X1 NAND2X1_814 (.gnd(gnd), .A(regs_2__9_), .Y(_4480_), .vdd(vdd), .B(raddr2_0_bF_buf96_), );
  NAND2X1 NAND2X1_815 (.gnd(gnd), .A(_4038__bF_buf7), .Y(_4481_), .vdd(vdd), .B(_4480_), );
  OAI21X1 OAI21X1_1743 (.gnd(gnd), .A(_4481_), .Y(_4482_), .vdd(vdd), .B(_4479_), .C(raddr2_2_bF_buf2_), );
  OAI22X1 OAI22X1_69 (.gnd(gnd), .A(_4478_), .Y(_4483_), .vdd(vdd), .B(_4482_), .C(_4476_), .D(_4473_), );
  NAND2X1 NAND2X1_816 (.gnd(gnd), .A(regs_10__9_), .Y(_4484_), .vdd(vdd), .B(raddr2_0_bF_buf95_), );
  OAI21X1 OAI21X1_1744 (.gnd(gnd), .A(_1920_), .Y(_4485_), .vdd(vdd), .B(raddr2_0_bF_buf94_), .C(_4484_), );
  NAND2X1 NAND2X1_817 (.gnd(gnd), .A(regs_8__9_), .Y(_4486_), .vdd(vdd), .B(raddr2_0_bF_buf93_), );
  OAI21X1 OAI21X1_1745 (.gnd(gnd), .A(_2018_), .Y(_4487_), .vdd(vdd), .B(raddr2_0_bF_buf92_), .C(_4486_), );
  MUX2X1 MUX2X1_387 (.gnd(gnd), .A(_4487_), .Y(_4488_), .vdd(vdd), .B(_4485_), .S(raddr2_1_bF_buf13_bF_buf2_), );
  NAND2X1 NAND2X1_818 (.gnd(gnd), .A(regs_14__9_), .Y(_4489_), .vdd(vdd), .B(raddr2_0_bF_buf91_), );
  OAI21X1 OAI21X1_1746 (.gnd(gnd), .A(_1723_), .Y(_4490_), .vdd(vdd), .B(raddr2_0_bF_buf90_), .C(_4489_), );
  NAND2X1 NAND2X1_819 (.gnd(gnd), .A(regs_12__9_), .Y(_4491_), .vdd(vdd), .B(raddr2_0_bF_buf89_), );
  OAI21X1 OAI21X1_1747 (.gnd(gnd), .A(_1821_), .Y(_4492_), .vdd(vdd), .B(raddr2_0_bF_buf88_), .C(_4491_), );
  MUX2X1 MUX2X1_388 (.gnd(gnd), .A(_4492_), .Y(_4493_), .vdd(vdd), .B(_4490_), .S(raddr2_1_bF_buf12_bF_buf2_), );
  MUX2X1 MUX2X1_389 (.gnd(gnd), .A(_4493_), .Y(_4494_), .vdd(vdd), .B(_4488_), .S(_4036__bF_buf8), );
  MUX2X1 MUX2X1_390 (.gnd(gnd), .A(_4494_), .Y(_4495_), .vdd(vdd), .B(_4483_), .S(_4033__bF_buf0), );
  MUX2X1 MUX2X1_391 (.gnd(gnd), .A(_4495_), .Y(_5512__9_), .vdd(vdd), .B(_4471_), .S(raddr2_4_bF_buf0_), );
  OAI21X1 OAI21X1_1748 (.gnd(gnd), .A(_2935_), .Y(_4496_), .vdd(vdd), .B(raddr2_0_bF_buf87_), .C(raddr2_1_bF_buf11_), );
  AOI21X1 AOI21X1_284 (.gnd(gnd), .A(regs_4__10_), .Y(_4497_), .vdd(vdd), .B(raddr2_0_bF_buf86_), .C(_4496_), );
  AND2X2 AND2X2_55 (.gnd(gnd), .A(regs_6__10_), .Y(_4498_), .vdd(vdd), .B(raddr2_0_bF_buf85_), );
  OAI21X1 OAI21X1_1749 (.gnd(gnd), .A(_2121_), .Y(_4499_), .vdd(vdd), .B(raddr2_0_bF_buf84_), .C(_4038__bF_buf6), );
  OAI21X1 OAI21X1_1750 (.gnd(gnd), .A(_4499_), .Y(_4500_), .vdd(vdd), .B(_4498_), .C(_4036__bF_buf7), );
  OAI21X1 OAI21X1_1751 (.gnd(gnd), .A(_2941_), .Y(_4501_), .vdd(vdd), .B(raddr2_0_bF_buf83_), .C(raddr2_1_bF_buf10_), );
  AOI21X1 AOI21X1_285 (.gnd(gnd), .A(regs_0__10_), .Y(_4502_), .vdd(vdd), .B(raddr2_0_bF_buf82_), .C(_4501_), );
  NOR2X1 NOR2X1_211 (.gnd(gnd), .A(raddr2_0_bF_buf81_), .Y(_4503_), .vdd(vdd), .B(_2944_), );
  NAND2X1 NAND2X1_820 (.gnd(gnd), .A(regs_2__10_), .Y(_4504_), .vdd(vdd), .B(raddr2_0_bF_buf80_), );
  NAND2X1 NAND2X1_821 (.gnd(gnd), .A(_4038__bF_buf5), .Y(_4505_), .vdd(vdd), .B(_4504_), );
  OAI21X1 OAI21X1_1752 (.gnd(gnd), .A(_4505_), .Y(_4506_), .vdd(vdd), .B(_4503_), .C(raddr2_2_bF_buf1_), );
  OAI22X1 OAI22X1_70 (.gnd(gnd), .A(_4502_), .Y(_4507_), .vdd(vdd), .B(_4506_), .C(_4500_), .D(_4497_), );
  NAND2X1 NAND2X1_822 (.gnd(gnd), .A(regs_10__10_), .Y(_4508_), .vdd(vdd), .B(raddr2_0_bF_buf79_), );
  OAI21X1 OAI21X1_1753 (.gnd(gnd), .A(_1922_), .Y(_4509_), .vdd(vdd), .B(raddr2_0_bF_buf78_), .C(_4508_), );
  NAND2X1 NAND2X1_823 (.gnd(gnd), .A(regs_8__10_), .Y(_4510_), .vdd(vdd), .B(raddr2_0_bF_buf77_), );
  OAI21X1 OAI21X1_1754 (.gnd(gnd), .A(_2020_), .Y(_4511_), .vdd(vdd), .B(raddr2_0_bF_buf76_), .C(_4510_), );
  MUX2X1 MUX2X1_392 (.gnd(gnd), .A(_4511_), .Y(_4512_), .vdd(vdd), .B(_4509_), .S(raddr2_1_bF_buf9_), );
  NAND2X1 NAND2X1_824 (.gnd(gnd), .A(regs_14__10_), .Y(_4513_), .vdd(vdd), .B(raddr2_0_bF_buf75_), );
  OAI21X1 OAI21X1_1755 (.gnd(gnd), .A(_1725_), .Y(_4514_), .vdd(vdd), .B(raddr2_0_bF_buf74_), .C(_4513_), );
  NAND2X1 NAND2X1_825 (.gnd(gnd), .A(regs_12__10_), .Y(_4515_), .vdd(vdd), .B(raddr2_0_bF_buf73_), );
  OAI21X1 OAI21X1_1756 (.gnd(gnd), .A(_1823_), .Y(_4516_), .vdd(vdd), .B(raddr2_0_bF_buf72_), .C(_4515_), );
  MUX2X1 MUX2X1_393 (.gnd(gnd), .A(_4516_), .Y(_4517_), .vdd(vdd), .B(_4514_), .S(raddr2_1_bF_buf8_), );
  MUX2X1 MUX2X1_394 (.gnd(gnd), .A(_4517_), .Y(_4518_), .vdd(vdd), .B(_4512_), .S(_4036__bF_buf6), );
  MUX2X1 MUX2X1_395 (.gnd(gnd), .A(_4518_), .Y(_4519_), .vdd(vdd), .B(_4507_), .S(_4033__bF_buf7), );
  OAI21X1 OAI21X1_1757 (.gnd(gnd), .A(_1625_), .Y(_4520_), .vdd(vdd), .B(raddr2_0_bF_buf71_), .C(raddr2_1_bF_buf7_), );
  AOI21X1 AOI21X1_286 (.gnd(gnd), .A(regs_16__10_), .Y(_4521_), .vdd(vdd), .B(raddr2_0_bF_buf70_), .C(_4520_), );
  NOR2X1 NOR2X1_212 (.gnd(gnd), .A(raddr2_0_bF_buf69_), .Y(_4522_), .vdd(vdd), .B(_1527_), );
  NAND2X1 NAND2X1_826 (.gnd(gnd), .A(regs_18__10_), .Y(_4523_), .vdd(vdd), .B(raddr2_0_bF_buf68_), );
  NAND2X1 NAND2X1_827 (.gnd(gnd), .A(_4038__bF_buf4), .Y(_4524_), .vdd(vdd), .B(_4523_), );
  OAI21X1 OAI21X1_1758 (.gnd(gnd), .A(_4524_), .Y(_4525_), .vdd(vdd), .B(_4522_), .C(raddr2_2_bF_buf0_), );
  OAI21X1 OAI21X1_1759 (.gnd(gnd), .A(_1428_), .Y(_4526_), .vdd(vdd), .B(raddr2_0_bF_buf67_), .C(raddr2_1_bF_buf6_), );
  AOI21X1 AOI21X1_287 (.gnd(gnd), .A(regs_20__10_), .Y(_4527_), .vdd(vdd), .B(raddr2_0_bF_buf66_), .C(_4526_), );
  AND2X2 AND2X2_56 (.gnd(gnd), .A(regs_22__10_), .Y(_4528_), .vdd(vdd), .B(raddr2_0_bF_buf65_), );
  OAI21X1 OAI21X1_1760 (.gnd(gnd), .A(_1330_), .Y(_4529_), .vdd(vdd), .B(raddr2_0_bF_buf64_), .C(_4038__bF_buf3), );
  OAI21X1 OAI21X1_1761 (.gnd(gnd), .A(_4529_), .Y(_4530_), .vdd(vdd), .B(_4528_), .C(_4036__bF_buf5), );
  OAI22X1 OAI22X1_71 (.gnd(gnd), .A(_4521_), .Y(_4531_), .vdd(vdd), .B(_4525_), .C(_4530_), .D(_4527_), );
  NAND2X1 NAND2X1_828 (.gnd(gnd), .A(regs_28__10_), .Y(_4532_), .vdd(vdd), .B(raddr2_0_bF_buf63_), );
  OAI21X1 OAI21X1_1762 (.gnd(gnd), .A(_2928_), .Y(_4533_), .vdd(vdd), .B(raddr2_0_bF_buf62_), .C(_4532_), );
  MUX2X1 MUX2X1_396 (.gnd(gnd), .A(_4533_), .Y(_4534_), .vdd(vdd), .B(regs_30__10_), .S(raddr2_1_bF_buf5_), );
  NAND2X1 NAND2X1_829 (.gnd(gnd), .A(regs_26__10_), .Y(_4535_), .vdd(vdd), .B(raddr2_0_bF_buf61_), );
  OAI21X1 OAI21X1_1763 (.gnd(gnd), .A(_1163_), .Y(_4536_), .vdd(vdd), .B(raddr2_0_bF_buf60_), .C(_4535_), );
  NAND2X1 NAND2X1_830 (.gnd(gnd), .A(regs_24__10_), .Y(_4537_), .vdd(vdd), .B(raddr2_0_bF_buf59_), );
  OAI21X1 OAI21X1_1764 (.gnd(gnd), .A(_2925_), .Y(_4538_), .vdd(vdd), .B(raddr2_0_bF_buf58_), .C(_4537_), );
  MUX2X1 MUX2X1_397 (.gnd(gnd), .A(_4538_), .Y(_4539_), .vdd(vdd), .B(_4536_), .S(raddr2_1_bF_buf4_), );
  MUX2X1 MUX2X1_398 (.gnd(gnd), .A(_4539_), .Y(_4540_), .vdd(vdd), .B(_4534_), .S(raddr2_2_bF_buf10_), );
  MUX2X1 MUX2X1_399 (.gnd(gnd), .A(_4540_), .Y(_4541_), .vdd(vdd), .B(_4531_), .S(_4033__bF_buf6), );
  MUX2X1 MUX2X1_400 (.gnd(gnd), .A(_4519_), .Y(_5512__10_), .vdd(vdd), .B(_4541_), .S(raddr2_4_bF_buf4_), );
  OAI21X1 OAI21X1_1765 (.gnd(gnd), .A(_2962_), .Y(_4542_), .vdd(vdd), .B(raddr2_0_bF_buf57_), .C(raddr2_1_bF_buf3_), );
  AOI21X1 AOI21X1_288 (.gnd(gnd), .A(regs_4__11_), .Y(_4543_), .vdd(vdd), .B(raddr2_0_bF_buf56_), .C(_4542_), );
  AND2X2 AND2X2_57 (.gnd(gnd), .A(regs_6__11_), .Y(_4544_), .vdd(vdd), .B(raddr2_0_bF_buf55_), );
  OAI21X1 OAI21X1_1766 (.gnd(gnd), .A(_2123_), .Y(_4545_), .vdd(vdd), .B(raddr2_0_bF_buf54_), .C(_4038__bF_buf2), );
  OAI21X1 OAI21X1_1767 (.gnd(gnd), .A(_4545_), .Y(_4546_), .vdd(vdd), .B(_4544_), .C(_4036__bF_buf4), );
  OAI21X1 OAI21X1_1768 (.gnd(gnd), .A(_2968_), .Y(_4547_), .vdd(vdd), .B(raddr2_0_bF_buf53_), .C(raddr2_1_bF_buf2_), );
  AOI21X1 AOI21X1_289 (.gnd(gnd), .A(regs_0__11_), .Y(_4548_), .vdd(vdd), .B(raddr2_0_bF_buf52_), .C(_4547_), );
  NOR2X1 NOR2X1_213 (.gnd(gnd), .A(raddr2_0_bF_buf51_), .Y(_4549_), .vdd(vdd), .B(_2971_), );
  NAND2X1 NAND2X1_831 (.gnd(gnd), .A(regs_2__11_), .Y(_4550_), .vdd(vdd), .B(raddr2_0_bF_buf50_), );
  NAND2X1 NAND2X1_832 (.gnd(gnd), .A(_4038__bF_buf1), .Y(_4551_), .vdd(vdd), .B(_4550_), );
  OAI21X1 OAI21X1_1769 (.gnd(gnd), .A(_4551_), .Y(_4552_), .vdd(vdd), .B(_4549_), .C(raddr2_2_bF_buf9_), );
  OAI22X1 OAI22X1_72 (.gnd(gnd), .A(_4548_), .Y(_4553_), .vdd(vdd), .B(_4552_), .C(_4546_), .D(_4543_), );
  NAND2X1 NAND2X1_833 (.gnd(gnd), .A(regs_10__11_), .Y(_4554_), .vdd(vdd), .B(raddr2_0_bF_buf49_), );
  OAI21X1 OAI21X1_1770 (.gnd(gnd), .A(_1924_), .Y(_4555_), .vdd(vdd), .B(raddr2_0_bF_buf48_), .C(_4554_), );
  NAND2X1 NAND2X1_834 (.gnd(gnd), .A(regs_8__11_), .Y(_4556_), .vdd(vdd), .B(raddr2_0_bF_buf47_), );
  OAI21X1 OAI21X1_1771 (.gnd(gnd), .A(_2022_), .Y(_4557_), .vdd(vdd), .B(raddr2_0_bF_buf46_), .C(_4556_), );
  MUX2X1 MUX2X1_401 (.gnd(gnd), .A(_4557_), .Y(_4558_), .vdd(vdd), .B(_4555_), .S(raddr2_1_bF_buf1_), );
  NAND2X1 NAND2X1_835 (.gnd(gnd), .A(regs_14__11_), .Y(_4559_), .vdd(vdd), .B(raddr2_0_bF_buf45_), );
  OAI21X1 OAI21X1_1772 (.gnd(gnd), .A(_1727_), .Y(_4560_), .vdd(vdd), .B(raddr2_0_bF_buf44_), .C(_4559_), );
  NAND2X1 NAND2X1_836 (.gnd(gnd), .A(regs_12__11_), .Y(_4561_), .vdd(vdd), .B(raddr2_0_bF_buf43_), );
  OAI21X1 OAI21X1_1773 (.gnd(gnd), .A(_1825_), .Y(_4562_), .vdd(vdd), .B(raddr2_0_bF_buf42_), .C(_4561_), );
  MUX2X1 MUX2X1_402 (.gnd(gnd), .A(_4562_), .Y(_4563_), .vdd(vdd), .B(_4560_), .S(raddr2_1_bF_buf0_), );
  MUX2X1 MUX2X1_403 (.gnd(gnd), .A(_4563_), .Y(_4564_), .vdd(vdd), .B(_4558_), .S(_4036__bF_buf3), );
  MUX2X1 MUX2X1_404 (.gnd(gnd), .A(_4564_), .Y(_4565_), .vdd(vdd), .B(_4553_), .S(_4033__bF_buf5), );
  OAI21X1 OAI21X1_1774 (.gnd(gnd), .A(_1627_), .Y(_4566_), .vdd(vdd), .B(raddr2_0_bF_buf41_), .C(raddr2_1_bF_buf14_bF_buf1_), );
  AOI21X1 AOI21X1_290 (.gnd(gnd), .A(regs_16__11_), .Y(_4567_), .vdd(vdd), .B(raddr2_0_bF_buf40_), .C(_4566_), );
  NOR2X1 NOR2X1_214 (.gnd(gnd), .A(raddr2_0_bF_buf39_), .Y(_4568_), .vdd(vdd), .B(_1529_), );
  NAND2X1 NAND2X1_837 (.gnd(gnd), .A(regs_18__11_), .Y(_4569_), .vdd(vdd), .B(raddr2_0_bF_buf38_), );
  NAND2X1 NAND2X1_838 (.gnd(gnd), .A(_4038__bF_buf0), .Y(_4570_), .vdd(vdd), .B(_4569_), );
  OAI21X1 OAI21X1_1775 (.gnd(gnd), .A(_4570_), .Y(_4571_), .vdd(vdd), .B(_4568_), .C(raddr2_2_bF_buf8_), );
  OAI21X1 OAI21X1_1776 (.gnd(gnd), .A(_1430_), .Y(_4572_), .vdd(vdd), .B(raddr2_0_bF_buf37_), .C(raddr2_1_bF_buf13_bF_buf1_), );
  AOI21X1 AOI21X1_291 (.gnd(gnd), .A(regs_20__11_), .Y(_4573_), .vdd(vdd), .B(raddr2_0_bF_buf36_), .C(_4572_), );
  AND2X2 AND2X2_58 (.gnd(gnd), .A(regs_22__11_), .Y(_4574_), .vdd(vdd), .B(raddr2_0_bF_buf35_), );
  OAI21X1 OAI21X1_1777 (.gnd(gnd), .A(_1332_), .Y(_4575_), .vdd(vdd), .B(raddr2_0_bF_buf34_), .C(_4038__bF_buf8), );
  OAI21X1 OAI21X1_1778 (.gnd(gnd), .A(_4575_), .Y(_4576_), .vdd(vdd), .B(_4574_), .C(_4036__bF_buf2), );
  OAI22X1 OAI22X1_73 (.gnd(gnd), .A(_4567_), .Y(_4577_), .vdd(vdd), .B(_4571_), .C(_4576_), .D(_4573_), );
  NAND2X1 NAND2X1_839 (.gnd(gnd), .A(regs_28__11_), .Y(_4578_), .vdd(vdd), .B(raddr2_0_bF_buf33_), );
  OAI21X1 OAI21X1_1779 (.gnd(gnd), .A(_3001_), .Y(_4579_), .vdd(vdd), .B(raddr2_0_bF_buf32_), .C(_4578_), );
  MUX2X1 MUX2X1_405 (.gnd(gnd), .A(_4579_), .Y(_4580_), .vdd(vdd), .B(regs_30__11_), .S(raddr2_1_bF_buf12_bF_buf1_), );
  NAND2X1 NAND2X1_840 (.gnd(gnd), .A(regs_26__11_), .Y(_4581_), .vdd(vdd), .B(raddr2_0_bF_buf31_), );
  OAI21X1 OAI21X1_1780 (.gnd(gnd), .A(_1165_), .Y(_4582_), .vdd(vdd), .B(raddr2_0_bF_buf30_), .C(_4581_), );
  NAND2X1 NAND2X1_841 (.gnd(gnd), .A(regs_24__11_), .Y(_4583_), .vdd(vdd), .B(raddr2_0_bF_buf29_), );
  OAI21X1 OAI21X1_1781 (.gnd(gnd), .A(_3007_), .Y(_4584_), .vdd(vdd), .B(raddr2_0_bF_buf28_), .C(_4583_), );
  MUX2X1 MUX2X1_406 (.gnd(gnd), .A(_4584_), .Y(_4585_), .vdd(vdd), .B(_4582_), .S(raddr2_1_bF_buf11_), );
  MUX2X1 MUX2X1_407 (.gnd(gnd), .A(_4585_), .Y(_4586_), .vdd(vdd), .B(_4580_), .S(raddr2_2_bF_buf7_), );
  MUX2X1 MUX2X1_408 (.gnd(gnd), .A(_4586_), .Y(_4587_), .vdd(vdd), .B(_4577_), .S(_4033__bF_buf4), );
  MUX2X1 MUX2X1_409 (.gnd(gnd), .A(_4565_), .Y(_5512__11_), .vdd(vdd), .B(_4587_), .S(raddr2_4_bF_buf3_), );
  OAI21X1 OAI21X1_1782 (.gnd(gnd), .A(_3013_), .Y(_4588_), .vdd(vdd), .B(raddr2_0_bF_buf27_), .C(raddr2_1_bF_buf10_), );
  AOI21X1 AOI21X1_292 (.gnd(gnd), .A(regs_4__12_), .Y(_4589_), .vdd(vdd), .B(raddr2_0_bF_buf26_), .C(_4588_), );
  AND2X2 AND2X2_59 (.gnd(gnd), .A(regs_6__12_), .Y(_4590_), .vdd(vdd), .B(raddr2_0_bF_buf25_), );
  OAI21X1 OAI21X1_1783 (.gnd(gnd), .A(_2125_), .Y(_4591_), .vdd(vdd), .B(raddr2_0_bF_buf24_), .C(_4038__bF_buf7), );
  OAI21X1 OAI21X1_1784 (.gnd(gnd), .A(_4591_), .Y(_4592_), .vdd(vdd), .B(_4590_), .C(_4036__bF_buf1), );
  OAI21X1 OAI21X1_1785 (.gnd(gnd), .A(_3019_), .Y(_4593_), .vdd(vdd), .B(raddr2_0_bF_buf23_), .C(raddr2_1_bF_buf9_), );
  AOI21X1 AOI21X1_293 (.gnd(gnd), .A(regs_0__12_), .Y(_4594_), .vdd(vdd), .B(raddr2_0_bF_buf22_), .C(_4593_), );
  NOR2X1 NOR2X1_215 (.gnd(gnd), .A(raddr2_0_bF_buf21_), .Y(_4595_), .vdd(vdd), .B(_3022_), );
  NAND2X1 NAND2X1_842 (.gnd(gnd), .A(regs_2__12_), .Y(_4596_), .vdd(vdd), .B(raddr2_0_bF_buf20_), );
  NAND2X1 NAND2X1_843 (.gnd(gnd), .A(_4038__bF_buf6), .Y(_4597_), .vdd(vdd), .B(_4596_), );
  OAI21X1 OAI21X1_1786 (.gnd(gnd), .A(_4597_), .Y(_4598_), .vdd(vdd), .B(_4595_), .C(raddr2_2_bF_buf6_), );
  OAI22X1 OAI22X1_74 (.gnd(gnd), .A(_4594_), .Y(_4599_), .vdd(vdd), .B(_4598_), .C(_4592_), .D(_4589_), );
  NAND2X1 NAND2X1_844 (.gnd(gnd), .A(regs_10__12_), .Y(_4600_), .vdd(vdd), .B(raddr2_0_bF_buf19_), );
  OAI21X1 OAI21X1_1787 (.gnd(gnd), .A(_1926_), .Y(_4601_), .vdd(vdd), .B(raddr2_0_bF_buf18_), .C(_4600_), );
  NAND2X1 NAND2X1_845 (.gnd(gnd), .A(regs_8__12_), .Y(_4602_), .vdd(vdd), .B(raddr2_0_bF_buf17_), );
  OAI21X1 OAI21X1_1788 (.gnd(gnd), .A(_2024_), .Y(_4603_), .vdd(vdd), .B(raddr2_0_bF_buf16_), .C(_4602_), );
  MUX2X1 MUX2X1_410 (.gnd(gnd), .A(_4603_), .Y(_4604_), .vdd(vdd), .B(_4601_), .S(raddr2_1_bF_buf8_), );
  NAND2X1 NAND2X1_846 (.gnd(gnd), .A(regs_14__12_), .Y(_4605_), .vdd(vdd), .B(raddr2_0_bF_buf15_), );
  OAI21X1 OAI21X1_1789 (.gnd(gnd), .A(_1729_), .Y(_4606_), .vdd(vdd), .B(raddr2_0_bF_buf14_), .C(_4605_), );
  NAND2X1 NAND2X1_847 (.gnd(gnd), .A(regs_12__12_), .Y(_4607_), .vdd(vdd), .B(raddr2_0_bF_buf13_), );
  OAI21X1 OAI21X1_1790 (.gnd(gnd), .A(_1827_), .Y(_4608_), .vdd(vdd), .B(raddr2_0_bF_buf12_), .C(_4607_), );
  MUX2X1 MUX2X1_411 (.gnd(gnd), .A(_4608_), .Y(_4609_), .vdd(vdd), .B(_4606_), .S(raddr2_1_bF_buf7_), );
  MUX2X1 MUX2X1_412 (.gnd(gnd), .A(_4609_), .Y(_4610_), .vdd(vdd), .B(_4604_), .S(_4036__bF_buf0), );
  MUX2X1 MUX2X1_413 (.gnd(gnd), .A(_4610_), .Y(_4611_), .vdd(vdd), .B(_4599_), .S(_4033__bF_buf3), );
  OAI21X1 OAI21X1_1791 (.gnd(gnd), .A(_1629_), .Y(_4612_), .vdd(vdd), .B(raddr2_0_bF_buf11_), .C(raddr2_1_bF_buf6_), );
  AOI21X1 AOI21X1_294 (.gnd(gnd), .A(regs_16__12_), .Y(_4613_), .vdd(vdd), .B(raddr2_0_bF_buf10_), .C(_4612_), );
  NOR2X1 NOR2X1_216 (.gnd(gnd), .A(raddr2_0_bF_buf9_), .Y(_4614_), .vdd(vdd), .B(_1531_), );
  NAND2X1 NAND2X1_848 (.gnd(gnd), .A(regs_18__12_), .Y(_4615_), .vdd(vdd), .B(raddr2_0_bF_buf8_), );
  NAND2X1 NAND2X1_849 (.gnd(gnd), .A(_4038__bF_buf5), .Y(_4616_), .vdd(vdd), .B(_4615_), );
  OAI21X1 OAI21X1_1792 (.gnd(gnd), .A(_4616_), .Y(_4617_), .vdd(vdd), .B(_4614_), .C(raddr2_2_bF_buf5_), );
  OAI21X1 OAI21X1_1793 (.gnd(gnd), .A(_1432_), .Y(_4618_), .vdd(vdd), .B(raddr2_0_bF_buf7_), .C(raddr2_1_bF_buf5_), );
  AOI21X1 AOI21X1_295 (.gnd(gnd), .A(regs_20__12_), .Y(_4619_), .vdd(vdd), .B(raddr2_0_bF_buf6_), .C(_4618_), );
  AND2X2 AND2X2_60 (.gnd(gnd), .A(regs_22__12_), .Y(_4620_), .vdd(vdd), .B(raddr2_0_bF_buf5_), );
  OAI21X1 OAI21X1_1794 (.gnd(gnd), .A(_1334_), .Y(_4621_), .vdd(vdd), .B(raddr2_0_bF_buf4_), .C(_4038__bF_buf4), );
  OAI21X1 OAI21X1_1795 (.gnd(gnd), .A(_4621_), .Y(_4622_), .vdd(vdd), .B(_4620_), .C(_4036__bF_buf8), );
  OAI22X1 OAI22X1_75 (.gnd(gnd), .A(_4613_), .Y(_4623_), .vdd(vdd), .B(_4617_), .C(_4622_), .D(_4619_), );
  NAND2X1 NAND2X1_850 (.gnd(gnd), .A(regs_28__12_), .Y(_4624_), .vdd(vdd), .B(raddr2_0_bF_buf3_), );
  OAI21X1 OAI21X1_1796 (.gnd(gnd), .A(_3052_), .Y(_4625_), .vdd(vdd), .B(raddr2_0_bF_buf2_), .C(_4624_), );
  MUX2X1 MUX2X1_414 (.gnd(gnd), .A(_4625_), .Y(_4626_), .vdd(vdd), .B(regs_30__12_), .S(raddr2_1_bF_buf4_), );
  NAND2X1 NAND2X1_851 (.gnd(gnd), .A(regs_26__12_), .Y(_4627_), .vdd(vdd), .B(raddr2_0_bF_buf1_), );
  OAI21X1 OAI21X1_1797 (.gnd(gnd), .A(_1167_), .Y(_4628_), .vdd(vdd), .B(raddr2_0_bF_buf0_), .C(_4627_), );
  NAND2X1 NAND2X1_852 (.gnd(gnd), .A(regs_24__12_), .Y(_4629_), .vdd(vdd), .B(raddr2_0_bF_buf96_), );
  OAI21X1 OAI21X1_1798 (.gnd(gnd), .A(_3058_), .Y(_4630_), .vdd(vdd), .B(raddr2_0_bF_buf95_), .C(_4629_), );
  MUX2X1 MUX2X1_415 (.gnd(gnd), .A(_4630_), .Y(_4631_), .vdd(vdd), .B(_4628_), .S(raddr2_1_bF_buf3_), );
  MUX2X1 MUX2X1_416 (.gnd(gnd), .A(_4631_), .Y(_4632_), .vdd(vdd), .B(_4626_), .S(raddr2_2_bF_buf4_), );
  MUX2X1 MUX2X1_417 (.gnd(gnd), .A(_4632_), .Y(_4633_), .vdd(vdd), .B(_4623_), .S(_4033__bF_buf2), );
  MUX2X1 MUX2X1_418 (.gnd(gnd), .A(_4611_), .Y(_5512__12_), .vdd(vdd), .B(_4633_), .S(raddr2_4_bF_buf2_), );
  OAI21X1 OAI21X1_1799 (.gnd(gnd), .A(_3064_), .Y(_4634_), .vdd(vdd), .B(raddr2_0_bF_buf94_), .C(raddr2_1_bF_buf2_), );
  AOI21X1 AOI21X1_296 (.gnd(gnd), .A(regs_4__13_), .Y(_4635_), .vdd(vdd), .B(raddr2_0_bF_buf93_), .C(_4634_), );
  AND2X2 AND2X2_61 (.gnd(gnd), .A(regs_6__13_), .Y(_4636_), .vdd(vdd), .B(raddr2_0_bF_buf92_), );
  OAI21X1 OAI21X1_1800 (.gnd(gnd), .A(_2127_), .Y(_4637_), .vdd(vdd), .B(raddr2_0_bF_buf91_), .C(_4038__bF_buf3), );
  OAI21X1 OAI21X1_1801 (.gnd(gnd), .A(_4637_), .Y(_4638_), .vdd(vdd), .B(_4636_), .C(_4036__bF_buf7), );
  OAI21X1 OAI21X1_1802 (.gnd(gnd), .A(_3070_), .Y(_4639_), .vdd(vdd), .B(raddr2_0_bF_buf90_), .C(raddr2_1_bF_buf1_), );
  AOI21X1 AOI21X1_297 (.gnd(gnd), .A(regs_0__13_), .Y(_4640_), .vdd(vdd), .B(raddr2_0_bF_buf89_), .C(_4639_), );
  NOR2X1 NOR2X1_217 (.gnd(gnd), .A(raddr2_0_bF_buf88_), .Y(_4641_), .vdd(vdd), .B(_3073_), );
  NAND2X1 NAND2X1_853 (.gnd(gnd), .A(regs_2__13_), .Y(_4642_), .vdd(vdd), .B(raddr2_0_bF_buf87_), );
  NAND2X1 NAND2X1_854 (.gnd(gnd), .A(_4038__bF_buf2), .Y(_4643_), .vdd(vdd), .B(_4642_), );
  OAI21X1 OAI21X1_1803 (.gnd(gnd), .A(_4643_), .Y(_4644_), .vdd(vdd), .B(_4641_), .C(raddr2_2_bF_buf3_), );
  OAI22X1 OAI22X1_76 (.gnd(gnd), .A(_4640_), .Y(_4645_), .vdd(vdd), .B(_4644_), .C(_4638_), .D(_4635_), );
  NAND2X1 NAND2X1_855 (.gnd(gnd), .A(regs_10__13_), .Y(_4646_), .vdd(vdd), .B(raddr2_0_bF_buf86_), );
  OAI21X1 OAI21X1_1804 (.gnd(gnd), .A(_1928_), .Y(_4647_), .vdd(vdd), .B(raddr2_0_bF_buf85_), .C(_4646_), );
  NAND2X1 NAND2X1_856 (.gnd(gnd), .A(regs_8__13_), .Y(_4648_), .vdd(vdd), .B(raddr2_0_bF_buf84_), );
  OAI21X1 OAI21X1_1805 (.gnd(gnd), .A(_2026_), .Y(_4649_), .vdd(vdd), .B(raddr2_0_bF_buf83_), .C(_4648_), );
  MUX2X1 MUX2X1_419 (.gnd(gnd), .A(_4649_), .Y(_4650_), .vdd(vdd), .B(_4647_), .S(raddr2_1_bF_buf0_), );
  NAND2X1 NAND2X1_857 (.gnd(gnd), .A(regs_14__13_), .Y(_4651_), .vdd(vdd), .B(raddr2_0_bF_buf82_), );
  OAI21X1 OAI21X1_1806 (.gnd(gnd), .A(_1731_), .Y(_4652_), .vdd(vdd), .B(raddr2_0_bF_buf81_), .C(_4651_), );
  NAND2X1 NAND2X1_858 (.gnd(gnd), .A(regs_12__13_), .Y(_4653_), .vdd(vdd), .B(raddr2_0_bF_buf80_), );
  OAI21X1 OAI21X1_1807 (.gnd(gnd), .A(_1829_), .Y(_4654_), .vdd(vdd), .B(raddr2_0_bF_buf79_), .C(_4653_), );
  MUX2X1 MUX2X1_420 (.gnd(gnd), .A(_4654_), .Y(_4655_), .vdd(vdd), .B(_4652_), .S(raddr2_1_bF_buf14_bF_buf0_), );
  MUX2X1 MUX2X1_421 (.gnd(gnd), .A(_4655_), .Y(_4656_), .vdd(vdd), .B(_4650_), .S(_4036__bF_buf6), );
  MUX2X1 MUX2X1_422 (.gnd(gnd), .A(_4656_), .Y(_4657_), .vdd(vdd), .B(_4645_), .S(_4033__bF_buf1), );
  OAI21X1 OAI21X1_1808 (.gnd(gnd), .A(_1631_), .Y(_4658_), .vdd(vdd), .B(raddr2_0_bF_buf78_), .C(raddr2_1_bF_buf13_bF_buf0_), );
  AOI21X1 AOI21X1_298 (.gnd(gnd), .A(regs_16__13_), .Y(_4659_), .vdd(vdd), .B(raddr2_0_bF_buf77_), .C(_4658_), );
  NOR2X1 NOR2X1_218 (.gnd(gnd), .A(raddr2_0_bF_buf76_), .Y(_4660_), .vdd(vdd), .B(_1533_), );
  NAND2X1 NAND2X1_859 (.gnd(gnd), .A(regs_18__13_), .Y(_4661_), .vdd(vdd), .B(raddr2_0_bF_buf75_), );
  NAND2X1 NAND2X1_860 (.gnd(gnd), .A(_4038__bF_buf1), .Y(_4662_), .vdd(vdd), .B(_4661_), );
  OAI21X1 OAI21X1_1809 (.gnd(gnd), .A(_4662_), .Y(_4663_), .vdd(vdd), .B(_4660_), .C(raddr2_2_bF_buf2_), );
  OAI21X1 OAI21X1_1810 (.gnd(gnd), .A(_1434_), .Y(_4664_), .vdd(vdd), .B(raddr2_0_bF_buf74_), .C(raddr2_1_bF_buf12_bF_buf0_), );
  AOI21X1 AOI21X1_299 (.gnd(gnd), .A(regs_20__13_), .Y(_4665_), .vdd(vdd), .B(raddr2_0_bF_buf73_), .C(_4664_), );
  AND2X2 AND2X2_62 (.gnd(gnd), .A(regs_22__13_), .Y(_4666_), .vdd(vdd), .B(raddr2_0_bF_buf72_), );
  OAI21X1 OAI21X1_1811 (.gnd(gnd), .A(_1336_), .Y(_4667_), .vdd(vdd), .B(raddr2_0_bF_buf71_), .C(_4038__bF_buf0), );
  OAI21X1 OAI21X1_1812 (.gnd(gnd), .A(_4667_), .Y(_4668_), .vdd(vdd), .B(_4666_), .C(_4036__bF_buf5), );
  OAI22X1 OAI22X1_77 (.gnd(gnd), .A(_4659_), .Y(_4669_), .vdd(vdd), .B(_4663_), .C(_4668_), .D(_4665_), );
  NAND2X1 NAND2X1_861 (.gnd(gnd), .A(regs_28__13_), .Y(_4670_), .vdd(vdd), .B(raddr2_0_bF_buf70_), );
  OAI21X1 OAI21X1_1813 (.gnd(gnd), .A(_3103_), .Y(_4671_), .vdd(vdd), .B(raddr2_0_bF_buf69_), .C(_4670_), );
  MUX2X1 MUX2X1_423 (.gnd(gnd), .A(_4671_), .Y(_4672_), .vdd(vdd), .B(regs_30__13_), .S(raddr2_1_bF_buf11_), );
  NAND2X1 NAND2X1_862 (.gnd(gnd), .A(regs_26__13_), .Y(_4673_), .vdd(vdd), .B(raddr2_0_bF_buf68_), );
  OAI21X1 OAI21X1_1814 (.gnd(gnd), .A(_1169_), .Y(_4674_), .vdd(vdd), .B(raddr2_0_bF_buf67_), .C(_4673_), );
  NAND2X1 NAND2X1_863 (.gnd(gnd), .A(regs_24__13_), .Y(_4675_), .vdd(vdd), .B(raddr2_0_bF_buf66_), );
  OAI21X1 OAI21X1_1815 (.gnd(gnd), .A(_3109_), .Y(_4676_), .vdd(vdd), .B(raddr2_0_bF_buf65_), .C(_4675_), );
  MUX2X1 MUX2X1_424 (.gnd(gnd), .A(_4676_), .Y(_4677_), .vdd(vdd), .B(_4674_), .S(raddr2_1_bF_buf10_), );
  MUX2X1 MUX2X1_425 (.gnd(gnd), .A(_4677_), .Y(_4678_), .vdd(vdd), .B(_4672_), .S(raddr2_2_bF_buf1_), );
  MUX2X1 MUX2X1_426 (.gnd(gnd), .A(_4678_), .Y(_4679_), .vdd(vdd), .B(_4669_), .S(_4033__bF_buf0), );
  MUX2X1 MUX2X1_427 (.gnd(gnd), .A(_4657_), .Y(_5512__13_), .vdd(vdd), .B(_4679_), .S(raddr2_4_bF_buf1_), );
  NAND2X1 NAND2X1_864 (.gnd(gnd), .A(regs_22__14_), .Y(_4680_), .vdd(vdd), .B(raddr2_0_bF_buf64_), );
  OAI21X1 OAI21X1_1816 (.gnd(gnd), .A(_1338_), .Y(_4681_), .vdd(vdd), .B(raddr2_0_bF_buf63_), .C(_4680_), );
  NAND2X1 NAND2X1_865 (.gnd(gnd), .A(regs_20__14_), .Y(_4682_), .vdd(vdd), .B(raddr2_0_bF_buf62_), );
  OAI21X1 OAI21X1_1817 (.gnd(gnd), .A(_1436_), .Y(_4683_), .vdd(vdd), .B(raddr2_0_bF_buf61_), .C(_4682_), );
  MUX2X1 MUX2X1_428 (.gnd(gnd), .A(_4683_), .Y(_4684_), .vdd(vdd), .B(_4681_), .S(raddr2_1_bF_buf9_), );
  NAND2X1 NAND2X1_866 (.gnd(gnd), .A(_4036__bF_buf4), .Y(_4685_), .vdd(vdd), .B(_4684_), );
  NAND2X1 NAND2X1_867 (.gnd(gnd), .A(regs_18__14_), .Y(_4686_), .vdd(vdd), .B(raddr2_0_bF_buf60_), );
  OAI21X1 OAI21X1_1818 (.gnd(gnd), .A(_1535_), .Y(_4687_), .vdd(vdd), .B(raddr2_0_bF_buf59_), .C(_4686_), );
  NAND2X1 NAND2X1_868 (.gnd(gnd), .A(regs_16__14_), .Y(_4688_), .vdd(vdd), .B(raddr2_0_bF_buf58_), );
  OAI21X1 OAI21X1_1819 (.gnd(gnd), .A(_1633_), .Y(_4689_), .vdd(vdd), .B(raddr2_0_bF_buf57_), .C(_4688_), );
  MUX2X1 MUX2X1_429 (.gnd(gnd), .A(_4689_), .Y(_4690_), .vdd(vdd), .B(_4687_), .S(raddr2_1_bF_buf8_), );
  AOI21X1 AOI21X1_300 (.gnd(gnd), .A(raddr2_2_bF_buf0_), .Y(_4691_), .vdd(vdd), .B(_4690_), .C(_4033__bF_buf7), );
  OAI21X1 OAI21X1_1820 (.gnd(gnd), .A(_1171_), .Y(_4692_), .vdd(vdd), .B(raddr2_0_bF_buf56_), .C(raddr2_2_bF_buf10_), );
  AOI21X1 AOI21X1_301 (.gnd(gnd), .A(regs_26__14_), .Y(_4693_), .vdd(vdd), .B(raddr2_0_bF_buf55_), .C(_4692_), );
  OAI21X1 OAI21X1_1821 (.gnd(gnd), .A(regs_30__14_), .Y(_4694_), .vdd(vdd), .B(raddr2_2_bF_buf9_), .C(_4038__bF_buf8), );
  OAI21X1 OAI21X1_1822 (.gnd(gnd), .A(_3130_), .Y(_4695_), .vdd(vdd), .B(raddr2_0_bF_buf54_), .C(raddr2_2_bF_buf8_), );
  AOI21X1 AOI21X1_302 (.gnd(gnd), .A(regs_24__14_), .Y(_4696_), .vdd(vdd), .B(raddr2_0_bF_buf53_), .C(_4695_), );
  NOR2X1 NOR2X1_219 (.gnd(gnd), .A(raddr2_0_bF_buf52_), .Y(_4697_), .vdd(vdd), .B(_3133_), );
  NAND2X1 NAND2X1_869 (.gnd(gnd), .A(regs_28__14_), .Y(_4698_), .vdd(vdd), .B(raddr2_0_bF_buf51_), );
  NAND2X1 NAND2X1_870 (.gnd(gnd), .A(_4036__bF_buf3), .Y(_4699_), .vdd(vdd), .B(_4698_), );
  OAI21X1 OAI21X1_1823 (.gnd(gnd), .A(_4699_), .Y(_4700_), .vdd(vdd), .B(_4697_), .C(raddr2_1_bF_buf7_), );
  OAI22X1 OAI22X1_78 (.gnd(gnd), .A(_4693_), .Y(_4701_), .vdd(vdd), .B(_4694_), .C(_4700_), .D(_4696_), );
  AOI22X1 AOI22X1_17 (.gnd(gnd), .A(_4701_), .Y(_4702_), .vdd(vdd), .B(_4033__bF_buf6), .C(_4685_), .D(_4691_), );
  OAI21X1 OAI21X1_1824 (.gnd(gnd), .A(_3140_), .Y(_4703_), .vdd(vdd), .B(raddr2_0_bF_buf50_), .C(raddr2_1_bF_buf6_), );
  AOI21X1 AOI21X1_303 (.gnd(gnd), .A(regs_4__14_), .Y(_4704_), .vdd(vdd), .B(raddr2_0_bF_buf49_), .C(_4703_), );
  AND2X2 AND2X2_63 (.gnd(gnd), .A(regs_6__14_), .Y(_4705_), .vdd(vdd), .B(raddr2_0_bF_buf48_), );
  OAI21X1 OAI21X1_1825 (.gnd(gnd), .A(_2129_), .Y(_4706_), .vdd(vdd), .B(raddr2_0_bF_buf47_), .C(_4038__bF_buf7), );
  OAI21X1 OAI21X1_1826 (.gnd(gnd), .A(_4706_), .Y(_4707_), .vdd(vdd), .B(_4705_), .C(_4036__bF_buf2), );
  OAI21X1 OAI21X1_1827 (.gnd(gnd), .A(_3146_), .Y(_4708_), .vdd(vdd), .B(raddr2_0_bF_buf46_), .C(raddr2_1_bF_buf5_), );
  AOI21X1 AOI21X1_304 (.gnd(gnd), .A(regs_0__14_), .Y(_4709_), .vdd(vdd), .B(raddr2_0_bF_buf45_), .C(_4708_), );
  NOR2X1 NOR2X1_220 (.gnd(gnd), .A(raddr2_0_bF_buf44_), .Y(_4710_), .vdd(vdd), .B(_3149_), );
  NAND2X1 NAND2X1_871 (.gnd(gnd), .A(regs_2__14_), .Y(_4711_), .vdd(vdd), .B(raddr2_0_bF_buf43_), );
  NAND2X1 NAND2X1_872 (.gnd(gnd), .A(_4038__bF_buf6), .Y(_4712_), .vdd(vdd), .B(_4711_), );
  OAI21X1 OAI21X1_1828 (.gnd(gnd), .A(_4712_), .Y(_4713_), .vdd(vdd), .B(_4710_), .C(raddr2_2_bF_buf7_), );
  OAI22X1 OAI22X1_79 (.gnd(gnd), .A(_4709_), .Y(_4714_), .vdd(vdd), .B(_4713_), .C(_4707_), .D(_4704_), );
  NAND2X1 NAND2X1_873 (.gnd(gnd), .A(regs_10__14_), .Y(_4715_), .vdd(vdd), .B(raddr2_0_bF_buf42_), );
  OAI21X1 OAI21X1_1829 (.gnd(gnd), .A(_1930_), .Y(_4716_), .vdd(vdd), .B(raddr2_0_bF_buf41_), .C(_4715_), );
  NAND2X1 NAND2X1_874 (.gnd(gnd), .A(regs_8__14_), .Y(_4717_), .vdd(vdd), .B(raddr2_0_bF_buf40_), );
  OAI21X1 OAI21X1_1830 (.gnd(gnd), .A(_2028_), .Y(_4718_), .vdd(vdd), .B(raddr2_0_bF_buf39_), .C(_4717_), );
  MUX2X1 MUX2X1_430 (.gnd(gnd), .A(_4718_), .Y(_4719_), .vdd(vdd), .B(_4716_), .S(raddr2_1_bF_buf4_), );
  NAND2X1 NAND2X1_875 (.gnd(gnd), .A(regs_14__14_), .Y(_4720_), .vdd(vdd), .B(raddr2_0_bF_buf38_), );
  OAI21X1 OAI21X1_1831 (.gnd(gnd), .A(_1733_), .Y(_4721_), .vdd(vdd), .B(raddr2_0_bF_buf37_), .C(_4720_), );
  NAND2X1 NAND2X1_876 (.gnd(gnd), .A(regs_12__14_), .Y(_4722_), .vdd(vdd), .B(raddr2_0_bF_buf36_), );
  OAI21X1 OAI21X1_1832 (.gnd(gnd), .A(_1831_), .Y(_4723_), .vdd(vdd), .B(raddr2_0_bF_buf35_), .C(_4722_), );
  MUX2X1 MUX2X1_431 (.gnd(gnd), .A(_4723_), .Y(_4724_), .vdd(vdd), .B(_4721_), .S(raddr2_1_bF_buf3_), );
  MUX2X1 MUX2X1_432 (.gnd(gnd), .A(_4724_), .Y(_4725_), .vdd(vdd), .B(_4719_), .S(_4036__bF_buf1), );
  MUX2X1 MUX2X1_433 (.gnd(gnd), .A(_4725_), .Y(_4726_), .vdd(vdd), .B(_4714_), .S(_4033__bF_buf5), );
  MUX2X1 MUX2X1_434 (.gnd(gnd), .A(_4726_), .Y(_5512__14_), .vdd(vdd), .B(_4702_), .S(raddr2_4_bF_buf0_), );
  NAND2X1 NAND2X1_877 (.gnd(gnd), .A(regs_22__15_), .Y(_4727_), .vdd(vdd), .B(raddr2_0_bF_buf34_), );
  OAI21X1 OAI21X1_1833 (.gnd(gnd), .A(_1340_), .Y(_4728_), .vdd(vdd), .B(raddr2_0_bF_buf33_), .C(_4727_), );
  NAND2X1 NAND2X1_878 (.gnd(gnd), .A(regs_20__15_), .Y(_4729_), .vdd(vdd), .B(raddr2_0_bF_buf32_), );
  OAI21X1 OAI21X1_1834 (.gnd(gnd), .A(_1438_), .Y(_4730_), .vdd(vdd), .B(raddr2_0_bF_buf31_), .C(_4729_), );
  MUX2X1 MUX2X1_435 (.gnd(gnd), .A(_4730_), .Y(_4731_), .vdd(vdd), .B(_4728_), .S(raddr2_1_bF_buf2_), );
  NAND2X1 NAND2X1_879 (.gnd(gnd), .A(_4036__bF_buf0), .Y(_4732_), .vdd(vdd), .B(_4731_), );
  NAND2X1 NAND2X1_880 (.gnd(gnd), .A(regs_18__15_), .Y(_4733_), .vdd(vdd), .B(raddr2_0_bF_buf30_), );
  OAI21X1 OAI21X1_1835 (.gnd(gnd), .A(_1537_), .Y(_4734_), .vdd(vdd), .B(raddr2_0_bF_buf29_), .C(_4733_), );
  NAND2X1 NAND2X1_881 (.gnd(gnd), .A(regs_16__15_), .Y(_4735_), .vdd(vdd), .B(raddr2_0_bF_buf28_), );
  OAI21X1 OAI21X1_1836 (.gnd(gnd), .A(_1635_), .Y(_4736_), .vdd(vdd), .B(raddr2_0_bF_buf27_), .C(_4735_), );
  MUX2X1 MUX2X1_436 (.gnd(gnd), .A(_4736_), .Y(_4737_), .vdd(vdd), .B(_4734_), .S(raddr2_1_bF_buf1_), );
  AOI21X1 AOI21X1_305 (.gnd(gnd), .A(raddr2_2_bF_buf6_), .Y(_4738_), .vdd(vdd), .B(_4737_), .C(_4033__bF_buf4), );
  OAI21X1 OAI21X1_1837 (.gnd(gnd), .A(_1173_), .Y(_4739_), .vdd(vdd), .B(raddr2_0_bF_buf26_), .C(raddr2_2_bF_buf5_), );
  AOI21X1 AOI21X1_306 (.gnd(gnd), .A(regs_26__15_), .Y(_4740_), .vdd(vdd), .B(raddr2_0_bF_buf25_), .C(_4739_), );
  OAI21X1 OAI21X1_1838 (.gnd(gnd), .A(regs_30__15_), .Y(_4741_), .vdd(vdd), .B(raddr2_2_bF_buf4_), .C(_4038__bF_buf5), );
  OAI21X1 OAI21X1_1839 (.gnd(gnd), .A(_3185_), .Y(_4742_), .vdd(vdd), .B(raddr2_0_bF_buf24_), .C(raddr2_2_bF_buf3_), );
  AOI21X1 AOI21X1_307 (.gnd(gnd), .A(regs_24__15_), .Y(_4743_), .vdd(vdd), .B(raddr2_0_bF_buf23_), .C(_4742_), );
  NOR2X1 NOR2X1_221 (.gnd(gnd), .A(raddr2_0_bF_buf22_), .Y(_4744_), .vdd(vdd), .B(_3179_), );
  NAND2X1 NAND2X1_882 (.gnd(gnd), .A(regs_28__15_), .Y(_4745_), .vdd(vdd), .B(raddr2_0_bF_buf21_), );
  NAND2X1 NAND2X1_883 (.gnd(gnd), .A(_4036__bF_buf8), .Y(_4746_), .vdd(vdd), .B(_4745_), );
  OAI21X1 OAI21X1_1840 (.gnd(gnd), .A(_4746_), .Y(_4747_), .vdd(vdd), .B(_4744_), .C(raddr2_1_bF_buf0_), );
  OAI22X1 OAI22X1_80 (.gnd(gnd), .A(_4740_), .Y(_4748_), .vdd(vdd), .B(_4741_), .C(_4747_), .D(_4743_), );
  AOI22X1 AOI22X1_18 (.gnd(gnd), .A(_4748_), .Y(_4749_), .vdd(vdd), .B(_4033__bF_buf3), .C(_4732_), .D(_4738_), );
  OAI21X1 OAI21X1_1841 (.gnd(gnd), .A(_3193_), .Y(_4750_), .vdd(vdd), .B(raddr2_0_bF_buf20_), .C(raddr2_1_bF_buf14_bF_buf3_), );
  AOI21X1 AOI21X1_308 (.gnd(gnd), .A(regs_4__15_), .Y(_4751_), .vdd(vdd), .B(raddr2_0_bF_buf19_), .C(_4750_), );
  AND2X2 AND2X2_64 (.gnd(gnd), .A(regs_6__15_), .Y(_4752_), .vdd(vdd), .B(raddr2_0_bF_buf18_), );
  OAI21X1 OAI21X1_1842 (.gnd(gnd), .A(_2131_), .Y(_4753_), .vdd(vdd), .B(raddr2_0_bF_buf17_), .C(_4038__bF_buf4), );
  OAI21X1 OAI21X1_1843 (.gnd(gnd), .A(_4753_), .Y(_4754_), .vdd(vdd), .B(_4752_), .C(_4036__bF_buf7), );
  OAI21X1 OAI21X1_1844 (.gnd(gnd), .A(_3200_), .Y(_4755_), .vdd(vdd), .B(raddr2_0_bF_buf16_), .C(raddr2_1_bF_buf13_bF_buf3_), );
  AOI21X1 AOI21X1_309 (.gnd(gnd), .A(regs_0__15_), .Y(_4756_), .vdd(vdd), .B(raddr2_0_bF_buf15_), .C(_4755_), );
  NOR2X1 NOR2X1_222 (.gnd(gnd), .A(raddr2_0_bF_buf14_), .Y(_4757_), .vdd(vdd), .B(_3197_), );
  NAND2X1 NAND2X1_884 (.gnd(gnd), .A(regs_2__15_), .Y(_4758_), .vdd(vdd), .B(raddr2_0_bF_buf13_), );
  NAND2X1 NAND2X1_885 (.gnd(gnd), .A(_4038__bF_buf3), .Y(_4759_), .vdd(vdd), .B(_4758_), );
  OAI21X1 OAI21X1_1845 (.gnd(gnd), .A(_4759_), .Y(_4760_), .vdd(vdd), .B(_4757_), .C(raddr2_2_bF_buf2_), );
  OAI22X1 OAI22X1_81 (.gnd(gnd), .A(_4756_), .Y(_4761_), .vdd(vdd), .B(_4760_), .C(_4754_), .D(_4751_), );
  NAND2X1 NAND2X1_886 (.gnd(gnd), .A(regs_10__15_), .Y(_4762_), .vdd(vdd), .B(raddr2_0_bF_buf12_), );
  OAI21X1 OAI21X1_1846 (.gnd(gnd), .A(_1932_), .Y(_4763_), .vdd(vdd), .B(raddr2_0_bF_buf11_), .C(_4762_), );
  NAND2X1 NAND2X1_887 (.gnd(gnd), .A(regs_8__15_), .Y(_4764_), .vdd(vdd), .B(raddr2_0_bF_buf10_), );
  OAI21X1 OAI21X1_1847 (.gnd(gnd), .A(_2030_), .Y(_4765_), .vdd(vdd), .B(raddr2_0_bF_buf9_), .C(_4764_), );
  MUX2X1 MUX2X1_437 (.gnd(gnd), .A(_4765_), .Y(_4766_), .vdd(vdd), .B(_4763_), .S(raddr2_1_bF_buf12_bF_buf3_), );
  NAND2X1 NAND2X1_888 (.gnd(gnd), .A(regs_14__15_), .Y(_4767_), .vdd(vdd), .B(raddr2_0_bF_buf8_), );
  OAI21X1 OAI21X1_1848 (.gnd(gnd), .A(_1735_), .Y(_4768_), .vdd(vdd), .B(raddr2_0_bF_buf7_), .C(_4767_), );
  NAND2X1 NAND2X1_889 (.gnd(gnd), .A(regs_12__15_), .Y(_4769_), .vdd(vdd), .B(raddr2_0_bF_buf6_), );
  OAI21X1 OAI21X1_1849 (.gnd(gnd), .A(_1833_), .Y(_4770_), .vdd(vdd), .B(raddr2_0_bF_buf5_), .C(_4769_), );
  MUX2X1 MUX2X1_438 (.gnd(gnd), .A(_4770_), .Y(_4771_), .vdd(vdd), .B(_4768_), .S(raddr2_1_bF_buf11_), );
  MUX2X1 MUX2X1_439 (.gnd(gnd), .A(_4771_), .Y(_4772_), .vdd(vdd), .B(_4766_), .S(_4036__bF_buf6), );
  MUX2X1 MUX2X1_440 (.gnd(gnd), .A(_4772_), .Y(_4773_), .vdd(vdd), .B(_4761_), .S(_4033__bF_buf2), );
  MUX2X1 MUX2X1_441 (.gnd(gnd), .A(_4773_), .Y(_5512__15_), .vdd(vdd), .B(_4749_), .S(raddr2_4_bF_buf4_), );
  NAND2X1 NAND2X1_890 (.gnd(gnd), .A(regs_22__16_), .Y(_4774_), .vdd(vdd), .B(raddr2_0_bF_buf4_), );
  OAI21X1 OAI21X1_1850 (.gnd(gnd), .A(_1342_), .Y(_4775_), .vdd(vdd), .B(raddr2_0_bF_buf3_), .C(_4774_), );
  NAND2X1 NAND2X1_891 (.gnd(gnd), .A(regs_20__16_), .Y(_4776_), .vdd(vdd), .B(raddr2_0_bF_buf2_), );
  OAI21X1 OAI21X1_1851 (.gnd(gnd), .A(_1440_), .Y(_4777_), .vdd(vdd), .B(raddr2_0_bF_buf1_), .C(_4776_), );
  MUX2X1 MUX2X1_442 (.gnd(gnd), .A(_4777_), .Y(_4778_), .vdd(vdd), .B(_4775_), .S(raddr2_1_bF_buf10_), );
  NAND2X1 NAND2X1_892 (.gnd(gnd), .A(_4036__bF_buf5), .Y(_4779_), .vdd(vdd), .B(_4778_), );
  NAND2X1 NAND2X1_893 (.gnd(gnd), .A(regs_18__16_), .Y(_4780_), .vdd(vdd), .B(raddr2_0_bF_buf0_), );
  OAI21X1 OAI21X1_1852 (.gnd(gnd), .A(_1539_), .Y(_4781_), .vdd(vdd), .B(raddr2_0_bF_buf96_), .C(_4780_), );
  NAND2X1 NAND2X1_894 (.gnd(gnd), .A(regs_16__16_), .Y(_4782_), .vdd(vdd), .B(raddr2_0_bF_buf95_), );
  OAI21X1 OAI21X1_1853 (.gnd(gnd), .A(_1637_), .Y(_4783_), .vdd(vdd), .B(raddr2_0_bF_buf94_), .C(_4782_), );
  MUX2X1 MUX2X1_443 (.gnd(gnd), .A(_4783_), .Y(_4784_), .vdd(vdd), .B(_4781_), .S(raddr2_1_bF_buf9_), );
  AOI21X1 AOI21X1_310 (.gnd(gnd), .A(raddr2_2_bF_buf1_), .Y(_4785_), .vdd(vdd), .B(_4784_), .C(_4033__bF_buf1), );
  OAI21X1 OAI21X1_1854 (.gnd(gnd), .A(_1175_), .Y(_4786_), .vdd(vdd), .B(raddr2_0_bF_buf93_), .C(raddr2_2_bF_buf0_), );
  AOI21X1 AOI21X1_311 (.gnd(gnd), .A(regs_26__16_), .Y(_4787_), .vdd(vdd), .B(raddr2_0_bF_buf92_), .C(_4786_), );
  OAI21X1 OAI21X1_1855 (.gnd(gnd), .A(regs_30__16_), .Y(_4788_), .vdd(vdd), .B(raddr2_2_bF_buf10_), .C(_4038__bF_buf2), );
  OAI21X1 OAI21X1_1856 (.gnd(gnd), .A(_3232_), .Y(_4789_), .vdd(vdd), .B(raddr2_0_bF_buf91_), .C(raddr2_2_bF_buf9_), );
  AOI21X1 AOI21X1_312 (.gnd(gnd), .A(regs_24__16_), .Y(_4790_), .vdd(vdd), .B(raddr2_0_bF_buf90_), .C(_4789_), );
  NOR2X1 NOR2X1_223 (.gnd(gnd), .A(raddr2_0_bF_buf89_), .Y(_4791_), .vdd(vdd), .B(_3235_), );
  NAND2X1 NAND2X1_895 (.gnd(gnd), .A(regs_28__16_), .Y(_4792_), .vdd(vdd), .B(raddr2_0_bF_buf88_), );
  NAND2X1 NAND2X1_896 (.gnd(gnd), .A(_4036__bF_buf4), .Y(_4793_), .vdd(vdd), .B(_4792_), );
  OAI21X1 OAI21X1_1857 (.gnd(gnd), .A(_4793_), .Y(_4794_), .vdd(vdd), .B(_4791_), .C(raddr2_1_bF_buf8_), );
  OAI22X1 OAI22X1_82 (.gnd(gnd), .A(_4787_), .Y(_4795_), .vdd(vdd), .B(_4788_), .C(_4794_), .D(_4790_), );
  AOI22X1 AOI22X1_19 (.gnd(gnd), .A(_4795_), .Y(_4796_), .vdd(vdd), .B(_4033__bF_buf0), .C(_4779_), .D(_4785_), );
  OAI21X1 OAI21X1_1858 (.gnd(gnd), .A(_3242_), .Y(_4797_), .vdd(vdd), .B(raddr2_0_bF_buf87_), .C(raddr2_1_bF_buf7_), );
  AOI21X1 AOI21X1_313 (.gnd(gnd), .A(regs_4__16_), .Y(_4798_), .vdd(vdd), .B(raddr2_0_bF_buf86_), .C(_4797_), );
  AND2X2 AND2X2_65 (.gnd(gnd), .A(regs_6__16_), .Y(_4799_), .vdd(vdd), .B(raddr2_0_bF_buf85_), );
  OAI21X1 OAI21X1_1859 (.gnd(gnd), .A(_2133_), .Y(_4800_), .vdd(vdd), .B(raddr2_0_bF_buf84_), .C(_4038__bF_buf1), );
  OAI21X1 OAI21X1_1860 (.gnd(gnd), .A(_4800_), .Y(_4801_), .vdd(vdd), .B(_4799_), .C(_4036__bF_buf3), );
  OAI21X1 OAI21X1_1861 (.gnd(gnd), .A(_3248_), .Y(_4802_), .vdd(vdd), .B(raddr2_0_bF_buf83_), .C(raddr2_1_bF_buf6_), );
  AOI21X1 AOI21X1_314 (.gnd(gnd), .A(regs_0__16_), .Y(_4803_), .vdd(vdd), .B(raddr2_0_bF_buf82_), .C(_4802_), );
  NOR2X1 NOR2X1_224 (.gnd(gnd), .A(raddr2_0_bF_buf81_), .Y(_4804_), .vdd(vdd), .B(_3251_), );
  NAND2X1 NAND2X1_897 (.gnd(gnd), .A(regs_2__16_), .Y(_4805_), .vdd(vdd), .B(raddr2_0_bF_buf80_), );
  NAND2X1 NAND2X1_898 (.gnd(gnd), .A(_4038__bF_buf0), .Y(_4806_), .vdd(vdd), .B(_4805_), );
  OAI21X1 OAI21X1_1862 (.gnd(gnd), .A(_4806_), .Y(_4807_), .vdd(vdd), .B(_4804_), .C(raddr2_2_bF_buf8_), );
  OAI22X1 OAI22X1_83 (.gnd(gnd), .A(_4803_), .Y(_4808_), .vdd(vdd), .B(_4807_), .C(_4801_), .D(_4798_), );
  NAND2X1 NAND2X1_899 (.gnd(gnd), .A(regs_10__16_), .Y(_4809_), .vdd(vdd), .B(raddr2_0_bF_buf79_), );
  OAI21X1 OAI21X1_1863 (.gnd(gnd), .A(_1934_), .Y(_4810_), .vdd(vdd), .B(raddr2_0_bF_buf78_), .C(_4809_), );
  NAND2X1 NAND2X1_900 (.gnd(gnd), .A(regs_8__16_), .Y(_4811_), .vdd(vdd), .B(raddr2_0_bF_buf77_), );
  OAI21X1 OAI21X1_1864 (.gnd(gnd), .A(_2032_), .Y(_4812_), .vdd(vdd), .B(raddr2_0_bF_buf76_), .C(_4811_), );
  MUX2X1 MUX2X1_444 (.gnd(gnd), .A(_4812_), .Y(_4813_), .vdd(vdd), .B(_4810_), .S(raddr2_1_bF_buf5_), );
  NAND2X1 NAND2X1_901 (.gnd(gnd), .A(regs_14__16_), .Y(_4814_), .vdd(vdd), .B(raddr2_0_bF_buf75_), );
  OAI21X1 OAI21X1_1865 (.gnd(gnd), .A(_1737_), .Y(_4815_), .vdd(vdd), .B(raddr2_0_bF_buf74_), .C(_4814_), );
  NAND2X1 NAND2X1_902 (.gnd(gnd), .A(regs_12__16_), .Y(_4816_), .vdd(vdd), .B(raddr2_0_bF_buf73_), );
  OAI21X1 OAI21X1_1866 (.gnd(gnd), .A(_1835_), .Y(_4817_), .vdd(vdd), .B(raddr2_0_bF_buf72_), .C(_4816_), );
  MUX2X1 MUX2X1_445 (.gnd(gnd), .A(_4817_), .Y(_4818_), .vdd(vdd), .B(_4815_), .S(raddr2_1_bF_buf4_), );
  MUX2X1 MUX2X1_446 (.gnd(gnd), .A(_4818_), .Y(_4819_), .vdd(vdd), .B(_4813_), .S(_4036__bF_buf2), );
  MUX2X1 MUX2X1_447 (.gnd(gnd), .A(_4819_), .Y(_4820_), .vdd(vdd), .B(_4808_), .S(_4033__bF_buf7), );
  MUX2X1 MUX2X1_448 (.gnd(gnd), .A(_4820_), .Y(_5512__16_), .vdd(vdd), .B(_4796_), .S(raddr2_4_bF_buf3_), );
  OAI21X1 OAI21X1_1867 (.gnd(gnd), .A(_1442_), .Y(_4821_), .vdd(vdd), .B(raddr2_0_bF_buf71_), .C(raddr2_1_bF_buf3_), );
  AOI21X1 AOI21X1_315 (.gnd(gnd), .A(regs_20__17_), .Y(_4822_), .vdd(vdd), .B(raddr2_0_bF_buf70_), .C(_4821_), );
  AND2X2 AND2X2_66 (.gnd(gnd), .A(regs_22__17_), .Y(_4823_), .vdd(vdd), .B(raddr2_0_bF_buf69_), );
  OAI21X1 OAI21X1_1868 (.gnd(gnd), .A(_1344_), .Y(_4824_), .vdd(vdd), .B(raddr2_0_bF_buf68_), .C(_4038__bF_buf8), );
  OAI21X1 OAI21X1_1869 (.gnd(gnd), .A(_4824_), .Y(_4825_), .vdd(vdd), .B(_4823_), .C(_4036__bF_buf1), );
  OAI21X1 OAI21X1_1870 (.gnd(gnd), .A(_1639_), .Y(_4826_), .vdd(vdd), .B(raddr2_0_bF_buf67_), .C(raddr2_1_bF_buf2_), );
  AOI21X1 AOI21X1_316 (.gnd(gnd), .A(regs_16__17_), .Y(_4827_), .vdd(vdd), .B(raddr2_0_bF_buf66_), .C(_4826_), );
  NOR2X1 NOR2X1_225 (.gnd(gnd), .A(raddr2_0_bF_buf65_), .Y(_4828_), .vdd(vdd), .B(_1541_), );
  NAND2X1 NAND2X1_903 (.gnd(gnd), .A(regs_18__17_), .Y(_4829_), .vdd(vdd), .B(raddr2_0_bF_buf64_), );
  NAND2X1 NAND2X1_904 (.gnd(gnd), .A(_4038__bF_buf7), .Y(_4830_), .vdd(vdd), .B(_4829_), );
  OAI21X1 OAI21X1_1871 (.gnd(gnd), .A(_4830_), .Y(_4831_), .vdd(vdd), .B(_4828_), .C(raddr2_2_bF_buf7_), );
  OAI22X1 OAI22X1_84 (.gnd(gnd), .A(_4827_), .Y(_4832_), .vdd(vdd), .B(_4831_), .C(_4825_), .D(_4822_), );
  NAND2X1 NAND2X1_905 (.gnd(gnd), .A(regs_28__17_), .Y(_4833_), .vdd(vdd), .B(raddr2_0_bF_buf63_), );
  OAI21X1 OAI21X1_1872 (.gnd(gnd), .A(_3287_), .Y(_4834_), .vdd(vdd), .B(raddr2_0_bF_buf62_), .C(_4833_), );
  MUX2X1 MUX2X1_449 (.gnd(gnd), .A(_4834_), .Y(_4835_), .vdd(vdd), .B(regs_30__17_), .S(raddr2_1_bF_buf1_), );
  NAND2X1 NAND2X1_906 (.gnd(gnd), .A(regs_26__17_), .Y(_4836_), .vdd(vdd), .B(raddr2_0_bF_buf61_), );
  OAI21X1 OAI21X1_1873 (.gnd(gnd), .A(_1177_), .Y(_4837_), .vdd(vdd), .B(raddr2_0_bF_buf60_), .C(_4836_), );
  NAND2X1 NAND2X1_907 (.gnd(gnd), .A(regs_24__17_), .Y(_4838_), .vdd(vdd), .B(raddr2_0_bF_buf59_), );
  OAI21X1 OAI21X1_1874 (.gnd(gnd), .A(_3284_), .Y(_4839_), .vdd(vdd), .B(raddr2_0_bF_buf58_), .C(_4838_), );
  MUX2X1 MUX2X1_450 (.gnd(gnd), .A(_4839_), .Y(_4840_), .vdd(vdd), .B(_4837_), .S(raddr2_1_bF_buf0_), );
  MUX2X1 MUX2X1_451 (.gnd(gnd), .A(_4840_), .Y(_4841_), .vdd(vdd), .B(_4835_), .S(raddr2_2_bF_buf6_), );
  MUX2X1 MUX2X1_452 (.gnd(gnd), .A(_4841_), .Y(_4842_), .vdd(vdd), .B(_4832_), .S(_4033__bF_buf6), );
  NAND2X1 NAND2X1_908 (.gnd(gnd), .A(regs_6__17_), .Y(_4843_), .vdd(vdd), .B(raddr2_0_bF_buf57_), );
  OAI21X1 OAI21X1_1875 (.gnd(gnd), .A(_2135_), .Y(_4844_), .vdd(vdd), .B(raddr2_0_bF_buf56_), .C(_4843_), );
  NAND2X1 NAND2X1_909 (.gnd(gnd), .A(regs_4__17_), .Y(_4845_), .vdd(vdd), .B(raddr2_0_bF_buf55_), );
  OAI21X1 OAI21X1_1876 (.gnd(gnd), .A(_3294_), .Y(_4846_), .vdd(vdd), .B(raddr2_0_bF_buf54_), .C(_4845_), );
  MUX2X1 MUX2X1_453 (.gnd(gnd), .A(_4846_), .Y(_4847_), .vdd(vdd), .B(_4844_), .S(raddr2_1_bF_buf14_bF_buf2_), );
  NAND2X1 NAND2X1_910 (.gnd(gnd), .A(regs_2__17_), .Y(_4848_), .vdd(vdd), .B(raddr2_0_bF_buf53_), );
  OAI21X1 OAI21X1_1877 (.gnd(gnd), .A(_3303_), .Y(_4849_), .vdd(vdd), .B(raddr2_0_bF_buf52_), .C(_4848_), );
  NAND2X1 NAND2X1_911 (.gnd(gnd), .A(regs_0__17_), .Y(_4850_), .vdd(vdd), .B(raddr2_0_bF_buf51_), );
  OAI21X1 OAI21X1_1878 (.gnd(gnd), .A(_3300_), .Y(_4851_), .vdd(vdd), .B(raddr2_0_bF_buf50_), .C(_4850_), );
  MUX2X1 MUX2X1_454 (.gnd(gnd), .A(_4851_), .Y(_4852_), .vdd(vdd), .B(_4849_), .S(raddr2_1_bF_buf13_bF_buf2_), );
  MUX2X1 MUX2X1_455 (.gnd(gnd), .A(_4852_), .Y(_4853_), .vdd(vdd), .B(_4847_), .S(raddr2_2_bF_buf5_), );
  NAND2X1 NAND2X1_912 (.gnd(gnd), .A(regs_14__17_), .Y(_4854_), .vdd(vdd), .B(raddr2_0_bF_buf49_), );
  OAI21X1 OAI21X1_1879 (.gnd(gnd), .A(_1739_), .Y(_4855_), .vdd(vdd), .B(raddr2_0_bF_buf48_), .C(_4854_), );
  NAND2X1 NAND2X1_913 (.gnd(gnd), .A(regs_12__17_), .Y(_4856_), .vdd(vdd), .B(raddr2_0_bF_buf47_), );
  OAI21X1 OAI21X1_1880 (.gnd(gnd), .A(_1837_), .Y(_4857_), .vdd(vdd), .B(raddr2_0_bF_buf46_), .C(_4856_), );
  MUX2X1 MUX2X1_456 (.gnd(gnd), .A(_4857_), .Y(_4858_), .vdd(vdd), .B(_4855_), .S(raddr2_1_bF_buf12_bF_buf2_), );
  NAND2X1 NAND2X1_914 (.gnd(gnd), .A(regs_10__17_), .Y(_4859_), .vdd(vdd), .B(raddr2_0_bF_buf45_), );
  OAI21X1 OAI21X1_1881 (.gnd(gnd), .A(_1936_), .Y(_4860_), .vdd(vdd), .B(raddr2_0_bF_buf44_), .C(_4859_), );
  NAND2X1 NAND2X1_915 (.gnd(gnd), .A(regs_8__17_), .Y(_4861_), .vdd(vdd), .B(raddr2_0_bF_buf43_), );
  OAI21X1 OAI21X1_1882 (.gnd(gnd), .A(_2034_), .Y(_4862_), .vdd(vdd), .B(raddr2_0_bF_buf42_), .C(_4861_), );
  MUX2X1 MUX2X1_457 (.gnd(gnd), .A(_4862_), .Y(_4863_), .vdd(vdd), .B(_4860_), .S(raddr2_1_bF_buf11_), );
  MUX2X1 MUX2X1_458 (.gnd(gnd), .A(_4863_), .Y(_4864_), .vdd(vdd), .B(_4858_), .S(raddr2_2_bF_buf4_), );
  MUX2X1 MUX2X1_459 (.gnd(gnd), .A(_4864_), .Y(_4865_), .vdd(vdd), .B(_4853_), .S(_4033__bF_buf5), );
  MUX2X1 MUX2X1_460 (.gnd(gnd), .A(_4865_), .Y(_5512__17_), .vdd(vdd), .B(_4842_), .S(raddr2_4_bF_buf2_), );
  NAND2X1 NAND2X1_916 (.gnd(gnd), .A(regs_22__18_), .Y(_4866_), .vdd(vdd), .B(raddr2_0_bF_buf41_), );
  OAI21X1 OAI21X1_1883 (.gnd(gnd), .A(_1346_), .Y(_4867_), .vdd(vdd), .B(raddr2_0_bF_buf40_), .C(_4866_), );
  NAND2X1 NAND2X1_917 (.gnd(gnd), .A(regs_20__18_), .Y(_4868_), .vdd(vdd), .B(raddr2_0_bF_buf39_), );
  OAI21X1 OAI21X1_1884 (.gnd(gnd), .A(_1444_), .Y(_4869_), .vdd(vdd), .B(raddr2_0_bF_buf38_), .C(_4868_), );
  MUX2X1 MUX2X1_461 (.gnd(gnd), .A(_4869_), .Y(_4870_), .vdd(vdd), .B(_4867_), .S(raddr2_1_bF_buf10_), );
  NAND2X1 NAND2X1_918 (.gnd(gnd), .A(_4036__bF_buf0), .Y(_4871_), .vdd(vdd), .B(_4870_), );
  NAND2X1 NAND2X1_919 (.gnd(gnd), .A(regs_18__18_), .Y(_4872_), .vdd(vdd), .B(raddr2_0_bF_buf37_), );
  OAI21X1 OAI21X1_1885 (.gnd(gnd), .A(_1543_), .Y(_4873_), .vdd(vdd), .B(raddr2_0_bF_buf36_), .C(_4872_), );
  NAND2X1 NAND2X1_920 (.gnd(gnd), .A(regs_16__18_), .Y(_4874_), .vdd(vdd), .B(raddr2_0_bF_buf35_), );
  OAI21X1 OAI21X1_1886 (.gnd(gnd), .A(_1641_), .Y(_4875_), .vdd(vdd), .B(raddr2_0_bF_buf34_), .C(_4874_), );
  MUX2X1 MUX2X1_462 (.gnd(gnd), .A(_4875_), .Y(_4876_), .vdd(vdd), .B(_4873_), .S(raddr2_1_bF_buf9_), );
  AOI21X1 AOI21X1_317 (.gnd(gnd), .A(raddr2_2_bF_buf3_), .Y(_4877_), .vdd(vdd), .B(_4876_), .C(_4033__bF_buf4), );
  OAI21X1 OAI21X1_1887 (.gnd(gnd), .A(_1179_), .Y(_4878_), .vdd(vdd), .B(raddr2_0_bF_buf33_), .C(raddr2_2_bF_buf2_), );
  AOI21X1 AOI21X1_318 (.gnd(gnd), .A(regs_26__18_), .Y(_4879_), .vdd(vdd), .B(raddr2_0_bF_buf32_), .C(_4878_), );
  OAI21X1 OAI21X1_1888 (.gnd(gnd), .A(regs_30__18_), .Y(_4880_), .vdd(vdd), .B(raddr2_2_bF_buf1_), .C(_4038__bF_buf6), );
  OAI21X1 OAI21X1_1889 (.gnd(gnd), .A(_3366_), .Y(_4881_), .vdd(vdd), .B(raddr2_0_bF_buf31_), .C(raddr2_2_bF_buf0_), );
  AOI21X1 AOI21X1_319 (.gnd(gnd), .A(regs_24__18_), .Y(_4882_), .vdd(vdd), .B(raddr2_0_bF_buf30_), .C(_4881_), );
  NOR2X1 NOR2X1_226 (.gnd(gnd), .A(raddr2_0_bF_buf29_), .Y(_4883_), .vdd(vdd), .B(_3360_), );
  NAND2X1 NAND2X1_921 (.gnd(gnd), .A(regs_28__18_), .Y(_4884_), .vdd(vdd), .B(raddr2_0_bF_buf28_), );
  NAND2X1 NAND2X1_922 (.gnd(gnd), .A(_4036__bF_buf8), .Y(_4885_), .vdd(vdd), .B(_4884_), );
  OAI21X1 OAI21X1_1890 (.gnd(gnd), .A(_4885_), .Y(_4886_), .vdd(vdd), .B(_4883_), .C(raddr2_1_bF_buf8_), );
  OAI22X1 OAI22X1_85 (.gnd(gnd), .A(_4879_), .Y(_4887_), .vdd(vdd), .B(_4880_), .C(_4886_), .D(_4882_), );
  AOI22X1 AOI22X1_20 (.gnd(gnd), .A(_4887_), .Y(_4888_), .vdd(vdd), .B(_4033__bF_buf3), .C(_4871_), .D(_4877_), );
  NAND2X1 NAND2X1_923 (.gnd(gnd), .A(regs_6__18_), .Y(_4889_), .vdd(vdd), .B(raddr2_0_bF_buf27_), );
  OAI21X1 OAI21X1_1891 (.gnd(gnd), .A(_2137_), .Y(_4890_), .vdd(vdd), .B(raddr2_0_bF_buf26_), .C(_4889_), );
  NAND2X1 NAND2X1_924 (.gnd(gnd), .A(regs_4__18_), .Y(_4891_), .vdd(vdd), .B(raddr2_0_bF_buf25_), );
  OAI21X1 OAI21X1_1892 (.gnd(gnd), .A(_3321_), .Y(_4892_), .vdd(vdd), .B(raddr2_0_bF_buf24_), .C(_4891_), );
  MUX2X1 MUX2X1_463 (.gnd(gnd), .A(_4892_), .Y(_4893_), .vdd(vdd), .B(_4890_), .S(raddr2_1_bF_buf7_), );
  NAND2X1 NAND2X1_925 (.gnd(gnd), .A(regs_2__18_), .Y(_4894_), .vdd(vdd), .B(raddr2_0_bF_buf23_), );
  OAI21X1 OAI21X1_1893 (.gnd(gnd), .A(_3330_), .Y(_4895_), .vdd(vdd), .B(raddr2_0_bF_buf22_), .C(_4894_), );
  NAND2X1 NAND2X1_926 (.gnd(gnd), .A(regs_0__18_), .Y(_4896_), .vdd(vdd), .B(raddr2_0_bF_buf21_), );
  OAI21X1 OAI21X1_1894 (.gnd(gnd), .A(_3327_), .Y(_4897_), .vdd(vdd), .B(raddr2_0_bF_buf20_), .C(_4896_), );
  MUX2X1 MUX2X1_464 (.gnd(gnd), .A(_4897_), .Y(_4898_), .vdd(vdd), .B(_4895_), .S(raddr2_1_bF_buf6_), );
  MUX2X1 MUX2X1_465 (.gnd(gnd), .A(_4898_), .Y(_4899_), .vdd(vdd), .B(_4893_), .S(raddr2_2_bF_buf10_), );
  NAND2X1 NAND2X1_927 (.gnd(gnd), .A(regs_10__18_), .Y(_4900_), .vdd(vdd), .B(raddr2_0_bF_buf19_), );
  OAI21X1 OAI21X1_1895 (.gnd(gnd), .A(_1938_), .Y(_4901_), .vdd(vdd), .B(raddr2_0_bF_buf18_), .C(_4900_), );
  NAND2X1 NAND2X1_928 (.gnd(gnd), .A(regs_8__18_), .Y(_4902_), .vdd(vdd), .B(raddr2_0_bF_buf17_), );
  OAI21X1 OAI21X1_1896 (.gnd(gnd), .A(_2036_), .Y(_4903_), .vdd(vdd), .B(raddr2_0_bF_buf16_), .C(_4902_), );
  MUX2X1 MUX2X1_466 (.gnd(gnd), .A(_4903_), .Y(_4904_), .vdd(vdd), .B(_4901_), .S(raddr2_1_bF_buf5_), );
  NAND2X1 NAND2X1_929 (.gnd(gnd), .A(regs_14__18_), .Y(_4905_), .vdd(vdd), .B(raddr2_0_bF_buf15_), );
  OAI21X1 OAI21X1_1897 (.gnd(gnd), .A(_1741_), .Y(_4906_), .vdd(vdd), .B(raddr2_0_bF_buf14_), .C(_4905_), );
  NAND2X1 NAND2X1_930 (.gnd(gnd), .A(regs_12__18_), .Y(_4907_), .vdd(vdd), .B(raddr2_0_bF_buf13_), );
  OAI21X1 OAI21X1_1898 (.gnd(gnd), .A(_1839_), .Y(_4908_), .vdd(vdd), .B(raddr2_0_bF_buf12_), .C(_4907_), );
  MUX2X1 MUX2X1_467 (.gnd(gnd), .A(_4908_), .Y(_4909_), .vdd(vdd), .B(_4906_), .S(raddr2_1_bF_buf4_), );
  MUX2X1 MUX2X1_468 (.gnd(gnd), .A(_4909_), .Y(_4910_), .vdd(vdd), .B(_4904_), .S(_4036__bF_buf7), );
  MUX2X1 MUX2X1_469 (.gnd(gnd), .A(_4910_), .Y(_4911_), .vdd(vdd), .B(_4899_), .S(_4033__bF_buf2), );
  MUX2X1 MUX2X1_470 (.gnd(gnd), .A(_4911_), .Y(_5512__18_), .vdd(vdd), .B(_4888_), .S(raddr2_4_bF_buf1_), );
  NAND2X1 NAND2X1_931 (.gnd(gnd), .A(regs_22__19_), .Y(_4912_), .vdd(vdd), .B(raddr2_0_bF_buf11_), );
  OAI21X1 OAI21X1_1899 (.gnd(gnd), .A(_1348_), .Y(_4913_), .vdd(vdd), .B(raddr2_0_bF_buf10_), .C(_4912_), );
  NAND2X1 NAND2X1_932 (.gnd(gnd), .A(regs_20__19_), .Y(_4914_), .vdd(vdd), .B(raddr2_0_bF_buf9_), );
  OAI21X1 OAI21X1_1900 (.gnd(gnd), .A(_1446_), .Y(_4915_), .vdd(vdd), .B(raddr2_0_bF_buf8_), .C(_4914_), );
  MUX2X1 MUX2X1_471 (.gnd(gnd), .A(_4915_), .Y(_4916_), .vdd(vdd), .B(_4913_), .S(raddr2_1_bF_buf3_), );
  NAND2X1 NAND2X1_933 (.gnd(gnd), .A(_4036__bF_buf6), .Y(_4917_), .vdd(vdd), .B(_4916_), );
  NAND2X1 NAND2X1_934 (.gnd(gnd), .A(regs_18__19_), .Y(_4918_), .vdd(vdd), .B(raddr2_0_bF_buf7_), );
  OAI21X1 OAI21X1_1901 (.gnd(gnd), .A(_1545_), .Y(_4919_), .vdd(vdd), .B(raddr2_0_bF_buf6_), .C(_4918_), );
  NAND2X1 NAND2X1_935 (.gnd(gnd), .A(regs_16__19_), .Y(_4920_), .vdd(vdd), .B(raddr2_0_bF_buf5_), );
  OAI21X1 OAI21X1_1902 (.gnd(gnd), .A(_1643_), .Y(_4921_), .vdd(vdd), .B(raddr2_0_bF_buf4_), .C(_4920_), );
  MUX2X1 MUX2X1_472 (.gnd(gnd), .A(_4921_), .Y(_4922_), .vdd(vdd), .B(_4919_), .S(raddr2_1_bF_buf2_), );
  AOI21X1 AOI21X1_320 (.gnd(gnd), .A(raddr2_2_bF_buf9_), .Y(_4923_), .vdd(vdd), .B(_4922_), .C(_4033__bF_buf1), );
  OAI21X1 OAI21X1_1903 (.gnd(gnd), .A(_1181_), .Y(_4924_), .vdd(vdd), .B(raddr2_0_bF_buf3_), .C(raddr2_2_bF_buf8_), );
  AOI21X1 AOI21X1_321 (.gnd(gnd), .A(regs_26__19_), .Y(_4925_), .vdd(vdd), .B(raddr2_0_bF_buf2_), .C(_4924_), );
  OAI21X1 OAI21X1_1904 (.gnd(gnd), .A(regs_30__19_), .Y(_4926_), .vdd(vdd), .B(raddr2_2_bF_buf7_), .C(_4038__bF_buf5), );
  OAI21X1 OAI21X1_1905 (.gnd(gnd), .A(_3387_), .Y(_4927_), .vdd(vdd), .B(raddr2_0_bF_buf1_), .C(raddr2_2_bF_buf6_), );
  AOI21X1 AOI21X1_322 (.gnd(gnd), .A(regs_24__19_), .Y(_4928_), .vdd(vdd), .B(raddr2_0_bF_buf0_), .C(_4927_), );
  NOR2X1 NOR2X1_227 (.gnd(gnd), .A(raddr2_0_bF_buf96_), .Y(_4929_), .vdd(vdd), .B(_3390_), );
  NAND2X1 NAND2X1_936 (.gnd(gnd), .A(regs_28__19_), .Y(_4930_), .vdd(vdd), .B(raddr2_0_bF_buf95_), );
  NAND2X1 NAND2X1_937 (.gnd(gnd), .A(_4036__bF_buf5), .Y(_4931_), .vdd(vdd), .B(_4930_), );
  OAI21X1 OAI21X1_1906 (.gnd(gnd), .A(_4931_), .Y(_4932_), .vdd(vdd), .B(_4929_), .C(raddr2_1_bF_buf1_), );
  OAI22X1 OAI22X1_86 (.gnd(gnd), .A(_4925_), .Y(_4933_), .vdd(vdd), .B(_4926_), .C(_4932_), .D(_4928_), );
  AOI22X1 AOI22X1_21 (.gnd(gnd), .A(_4933_), .Y(_4934_), .vdd(vdd), .B(_4033__bF_buf0), .C(_4917_), .D(_4923_), );
  NAND2X1 NAND2X1_938 (.gnd(gnd), .A(regs_6__19_), .Y(_4935_), .vdd(vdd), .B(raddr2_0_bF_buf94_), );
  OAI21X1 OAI21X1_1907 (.gnd(gnd), .A(_2139_), .Y(_4936_), .vdd(vdd), .B(raddr2_0_bF_buf93_), .C(_4935_), );
  NAND2X1 NAND2X1_939 (.gnd(gnd), .A(regs_4__19_), .Y(_4937_), .vdd(vdd), .B(raddr2_0_bF_buf92_), );
  OAI21X1 OAI21X1_1908 (.gnd(gnd), .A(_3399_), .Y(_4938_), .vdd(vdd), .B(raddr2_0_bF_buf91_), .C(_4937_), );
  MUX2X1 MUX2X1_473 (.gnd(gnd), .A(_4938_), .Y(_4939_), .vdd(vdd), .B(_4936_), .S(raddr2_1_bF_buf0_), );
  NAND2X1 NAND2X1_940 (.gnd(gnd), .A(regs_2__19_), .Y(_4940_), .vdd(vdd), .B(raddr2_0_bF_buf90_), );
  OAI21X1 OAI21X1_1909 (.gnd(gnd), .A(_3403_), .Y(_4941_), .vdd(vdd), .B(raddr2_0_bF_buf89_), .C(_4940_), );
  NAND2X1 NAND2X1_941 (.gnd(gnd), .A(regs_0__19_), .Y(_4942_), .vdd(vdd), .B(raddr2_0_bF_buf88_), );
  OAI21X1 OAI21X1_1910 (.gnd(gnd), .A(_3406_), .Y(_4943_), .vdd(vdd), .B(raddr2_0_bF_buf87_), .C(_4942_), );
  MUX2X1 MUX2X1_474 (.gnd(gnd), .A(_4943_), .Y(_4944_), .vdd(vdd), .B(_4941_), .S(raddr2_1_bF_buf14_bF_buf1_), );
  MUX2X1 MUX2X1_475 (.gnd(gnd), .A(_4944_), .Y(_4945_), .vdd(vdd), .B(_4939_), .S(raddr2_2_bF_buf5_), );
  NAND2X1 NAND2X1_942 (.gnd(gnd), .A(regs_10__19_), .Y(_4946_), .vdd(vdd), .B(raddr2_0_bF_buf86_), );
  OAI21X1 OAI21X1_1911 (.gnd(gnd), .A(_1940_), .Y(_4947_), .vdd(vdd), .B(raddr2_0_bF_buf85_), .C(_4946_), );
  NAND2X1 NAND2X1_943 (.gnd(gnd), .A(regs_8__19_), .Y(_4948_), .vdd(vdd), .B(raddr2_0_bF_buf84_), );
  OAI21X1 OAI21X1_1912 (.gnd(gnd), .A(_2038_), .Y(_4949_), .vdd(vdd), .B(raddr2_0_bF_buf83_), .C(_4948_), );
  MUX2X1 MUX2X1_476 (.gnd(gnd), .A(_4949_), .Y(_4950_), .vdd(vdd), .B(_4947_), .S(raddr2_1_bF_buf13_bF_buf1_), );
  NAND2X1 NAND2X1_944 (.gnd(gnd), .A(regs_14__19_), .Y(_4951_), .vdd(vdd), .B(raddr2_0_bF_buf82_), );
  OAI21X1 OAI21X1_1913 (.gnd(gnd), .A(_1743_), .Y(_4952_), .vdd(vdd), .B(raddr2_0_bF_buf81_), .C(_4951_), );
  NAND2X1 NAND2X1_945 (.gnd(gnd), .A(regs_12__19_), .Y(_4953_), .vdd(vdd), .B(raddr2_0_bF_buf80_), );
  OAI21X1 OAI21X1_1914 (.gnd(gnd), .A(_1841_), .Y(_4954_), .vdd(vdd), .B(raddr2_0_bF_buf79_), .C(_4953_), );
  MUX2X1 MUX2X1_477 (.gnd(gnd), .A(_4954_), .Y(_4955_), .vdd(vdd), .B(_4952_), .S(raddr2_1_bF_buf12_bF_buf1_), );
  MUX2X1 MUX2X1_478 (.gnd(gnd), .A(_4955_), .Y(_4956_), .vdd(vdd), .B(_4950_), .S(_4036__bF_buf4), );
  MUX2X1 MUX2X1_479 (.gnd(gnd), .A(_4956_), .Y(_4957_), .vdd(vdd), .B(_4945_), .S(_4033__bF_buf7), );
  MUX2X1 MUX2X1_480 (.gnd(gnd), .A(_4957_), .Y(_5512__19_), .vdd(vdd), .B(_4934_), .S(raddr2_4_bF_buf0_), );
  NAND2X1 NAND2X1_946 (.gnd(gnd), .A(regs_22__20_), .Y(_4958_), .vdd(vdd), .B(raddr2_0_bF_buf78_), );
  OAI21X1 OAI21X1_1915 (.gnd(gnd), .A(_1350_), .Y(_4959_), .vdd(vdd), .B(raddr2_0_bF_buf77_), .C(_4958_), );
  NAND2X1 NAND2X1_947 (.gnd(gnd), .A(regs_20__20_), .Y(_4960_), .vdd(vdd), .B(raddr2_0_bF_buf76_), );
  OAI21X1 OAI21X1_1916 (.gnd(gnd), .A(_1448_), .Y(_4961_), .vdd(vdd), .B(raddr2_0_bF_buf75_), .C(_4960_), );
  MUX2X1 MUX2X1_481 (.gnd(gnd), .A(_4961_), .Y(_4962_), .vdd(vdd), .B(_4959_), .S(raddr2_1_bF_buf11_), );
  NAND2X1 NAND2X1_948 (.gnd(gnd), .A(_4036__bF_buf3), .Y(_4963_), .vdd(vdd), .B(_4962_), );
  NAND2X1 NAND2X1_949 (.gnd(gnd), .A(regs_18__20_), .Y(_4964_), .vdd(vdd), .B(raddr2_0_bF_buf74_), );
  OAI21X1 OAI21X1_1917 (.gnd(gnd), .A(_1547_), .Y(_4965_), .vdd(vdd), .B(raddr2_0_bF_buf73_), .C(_4964_), );
  NAND2X1 NAND2X1_950 (.gnd(gnd), .A(regs_16__20_), .Y(_4966_), .vdd(vdd), .B(raddr2_0_bF_buf72_), );
  OAI21X1 OAI21X1_1918 (.gnd(gnd), .A(_1645_), .Y(_4967_), .vdd(vdd), .B(raddr2_0_bF_buf71_), .C(_4966_), );
  MUX2X1 MUX2X1_482 (.gnd(gnd), .A(_4967_), .Y(_4968_), .vdd(vdd), .B(_4965_), .S(raddr2_1_bF_buf10_), );
  AOI21X1 AOI21X1_323 (.gnd(gnd), .A(raddr2_2_bF_buf4_), .Y(_4969_), .vdd(vdd), .B(_4968_), .C(_4033__bF_buf6), );
  OAI21X1 OAI21X1_1919 (.gnd(gnd), .A(_1183_), .Y(_4970_), .vdd(vdd), .B(raddr2_0_bF_buf70_), .C(raddr2_2_bF_buf3_), );
  AOI21X1 AOI21X1_324 (.gnd(gnd), .A(regs_26__20_), .Y(_4971_), .vdd(vdd), .B(raddr2_0_bF_buf69_), .C(_4970_), );
  OAI21X1 OAI21X1_1920 (.gnd(gnd), .A(regs_30__20_), .Y(_4972_), .vdd(vdd), .B(raddr2_2_bF_buf2_), .C(_4038__bF_buf4), );
  OAI21X1 OAI21X1_1921 (.gnd(gnd), .A(_3468_), .Y(_4973_), .vdd(vdd), .B(raddr2_0_bF_buf68_), .C(raddr2_2_bF_buf1_), );
  AOI21X1 AOI21X1_325 (.gnd(gnd), .A(regs_24__20_), .Y(_4974_), .vdd(vdd), .B(raddr2_0_bF_buf67_), .C(_4973_), );
  NOR2X1 NOR2X1_228 (.gnd(gnd), .A(raddr2_0_bF_buf66_), .Y(_4975_), .vdd(vdd), .B(_3462_), );
  NAND2X1 NAND2X1_951 (.gnd(gnd), .A(regs_28__20_), .Y(_4976_), .vdd(vdd), .B(raddr2_0_bF_buf65_), );
  NAND2X1 NAND2X1_952 (.gnd(gnd), .A(_4036__bF_buf2), .Y(_4977_), .vdd(vdd), .B(_4976_), );
  OAI21X1 OAI21X1_1922 (.gnd(gnd), .A(_4977_), .Y(_4978_), .vdd(vdd), .B(_4975_), .C(raddr2_1_bF_buf9_), );
  OAI22X1 OAI22X1_87 (.gnd(gnd), .A(_4971_), .Y(_4979_), .vdd(vdd), .B(_4972_), .C(_4978_), .D(_4974_), );
  AOI22X1 AOI22X1_22 (.gnd(gnd), .A(_4979_), .Y(_4980_), .vdd(vdd), .B(_4033__bF_buf5), .C(_4963_), .D(_4969_), );
  NAND2X1 NAND2X1_953 (.gnd(gnd), .A(regs_6__20_), .Y(_4981_), .vdd(vdd), .B(raddr2_0_bF_buf64_), );
  OAI21X1 OAI21X1_1923 (.gnd(gnd), .A(_2141_), .Y(_4982_), .vdd(vdd), .B(raddr2_0_bF_buf63_), .C(_4981_), );
  NAND2X1 NAND2X1_954 (.gnd(gnd), .A(regs_4__20_), .Y(_4983_), .vdd(vdd), .B(raddr2_0_bF_buf62_), );
  OAI21X1 OAI21X1_1924 (.gnd(gnd), .A(_3423_), .Y(_4984_), .vdd(vdd), .B(raddr2_0_bF_buf61_), .C(_4983_), );
  MUX2X1 MUX2X1_483 (.gnd(gnd), .A(_4984_), .Y(_4985_), .vdd(vdd), .B(_4982_), .S(raddr2_1_bF_buf8_), );
  NAND2X1 NAND2X1_955 (.gnd(gnd), .A(regs_2__20_), .Y(_4986_), .vdd(vdd), .B(raddr2_0_bF_buf60_), );
  OAI21X1 OAI21X1_1925 (.gnd(gnd), .A(_3432_), .Y(_4987_), .vdd(vdd), .B(raddr2_0_bF_buf59_), .C(_4986_), );
  NAND2X1 NAND2X1_956 (.gnd(gnd), .A(regs_0__20_), .Y(_4988_), .vdd(vdd), .B(raddr2_0_bF_buf58_), );
  OAI21X1 OAI21X1_1926 (.gnd(gnd), .A(_3429_), .Y(_4989_), .vdd(vdd), .B(raddr2_0_bF_buf57_), .C(_4988_), );
  MUX2X1 MUX2X1_484 (.gnd(gnd), .A(_4989_), .Y(_4990_), .vdd(vdd), .B(_4987_), .S(raddr2_1_bF_buf7_), );
  MUX2X1 MUX2X1_485 (.gnd(gnd), .A(_4990_), .Y(_4991_), .vdd(vdd), .B(_4985_), .S(raddr2_2_bF_buf0_), );
  NAND2X1 NAND2X1_957 (.gnd(gnd), .A(regs_10__20_), .Y(_4992_), .vdd(vdd), .B(raddr2_0_bF_buf56_), );
  OAI21X1 OAI21X1_1927 (.gnd(gnd), .A(_1942_), .Y(_4993_), .vdd(vdd), .B(raddr2_0_bF_buf55_), .C(_4992_), );
  NAND2X1 NAND2X1_958 (.gnd(gnd), .A(regs_8__20_), .Y(_4994_), .vdd(vdd), .B(raddr2_0_bF_buf54_), );
  OAI21X1 OAI21X1_1928 (.gnd(gnd), .A(_2040_), .Y(_4995_), .vdd(vdd), .B(raddr2_0_bF_buf53_), .C(_4994_), );
  MUX2X1 MUX2X1_486 (.gnd(gnd), .A(_4995_), .Y(_4996_), .vdd(vdd), .B(_4993_), .S(raddr2_1_bF_buf6_), );
  NAND2X1 NAND2X1_959 (.gnd(gnd), .A(regs_14__20_), .Y(_4997_), .vdd(vdd), .B(raddr2_0_bF_buf52_), );
  OAI21X1 OAI21X1_1929 (.gnd(gnd), .A(_1745_), .Y(_4998_), .vdd(vdd), .B(raddr2_0_bF_buf51_), .C(_4997_), );
  NAND2X1 NAND2X1_960 (.gnd(gnd), .A(regs_12__20_), .Y(_4999_), .vdd(vdd), .B(raddr2_0_bF_buf50_), );
  OAI21X1 OAI21X1_1930 (.gnd(gnd), .A(_1843_), .Y(_5000_), .vdd(vdd), .B(raddr2_0_bF_buf49_), .C(_4999_), );
  MUX2X1 MUX2X1_487 (.gnd(gnd), .A(_5000_), .Y(_5001_), .vdd(vdd), .B(_4998_), .S(raddr2_1_bF_buf5_), );
  MUX2X1 MUX2X1_488 (.gnd(gnd), .A(_5001_), .Y(_5002_), .vdd(vdd), .B(_4996_), .S(_4036__bF_buf1), );
  MUX2X1 MUX2X1_489 (.gnd(gnd), .A(_5002_), .Y(_5003_), .vdd(vdd), .B(_4991_), .S(_4033__bF_buf4), );
  MUX2X1 MUX2X1_490 (.gnd(gnd), .A(_5003_), .Y(_5512__20_), .vdd(vdd), .B(_4980_), .S(raddr2_4_bF_buf4_), );
  OAI21X1 OAI21X1_1931 (.gnd(gnd), .A(_1450_), .Y(_5004_), .vdd(vdd), .B(raddr2_0_bF_buf48_), .C(raddr2_1_bF_buf4_), );
  AOI21X1 AOI21X1_326 (.gnd(gnd), .A(regs_20__21_), .Y(_5005_), .vdd(vdd), .B(raddr2_0_bF_buf47_), .C(_5004_), );
  AND2X2 AND2X2_67 (.gnd(gnd), .A(regs_22__21_), .Y(_5006_), .vdd(vdd), .B(raddr2_0_bF_buf46_), );
  OAI21X1 OAI21X1_1932 (.gnd(gnd), .A(_1352_), .Y(_5007_), .vdd(vdd), .B(raddr2_0_bF_buf45_), .C(_4038__bF_buf3), );
  OAI21X1 OAI21X1_1933 (.gnd(gnd), .A(_5007_), .Y(_5008_), .vdd(vdd), .B(_5006_), .C(_4036__bF_buf0), );
  OAI21X1 OAI21X1_1934 (.gnd(gnd), .A(_1647_), .Y(_5009_), .vdd(vdd), .B(raddr2_0_bF_buf44_), .C(raddr2_1_bF_buf3_), );
  AOI21X1 AOI21X1_327 (.gnd(gnd), .A(regs_16__21_), .Y(_5010_), .vdd(vdd), .B(raddr2_0_bF_buf43_), .C(_5009_), );
  NOR2X1 NOR2X1_229 (.gnd(gnd), .A(raddr2_0_bF_buf42_), .Y(_5011_), .vdd(vdd), .B(_1549_), );
  NAND2X1 NAND2X1_961 (.gnd(gnd), .A(regs_18__21_), .Y(_5012_), .vdd(vdd), .B(raddr2_0_bF_buf41_), );
  NAND2X1 NAND2X1_962 (.gnd(gnd), .A(_4038__bF_buf2), .Y(_5013_), .vdd(vdd), .B(_5012_), );
  OAI21X1 OAI21X1_1935 (.gnd(gnd), .A(_5013_), .Y(_5014_), .vdd(vdd), .B(_5011_), .C(raddr2_2_bF_buf10_), );
  OAI22X1 OAI22X1_88 (.gnd(gnd), .A(_5010_), .Y(_5015_), .vdd(vdd), .B(_5014_), .C(_5008_), .D(_5005_), );
  NAND2X1 NAND2X1_963 (.gnd(gnd), .A(regs_28__21_), .Y(_5016_), .vdd(vdd), .B(raddr2_0_bF_buf40_), );
  OAI21X1 OAI21X1_1936 (.gnd(gnd), .A(_3513_), .Y(_5017_), .vdd(vdd), .B(raddr2_0_bF_buf39_), .C(_5016_), );
  MUX2X1 MUX2X1_491 (.gnd(gnd), .A(_5017_), .Y(_5018_), .vdd(vdd), .B(regs_30__21_), .S(raddr2_1_bF_buf2_), );
  NAND2X1 NAND2X1_964 (.gnd(gnd), .A(regs_26__21_), .Y(_5019_), .vdd(vdd), .B(raddr2_0_bF_buf38_), );
  OAI21X1 OAI21X1_1937 (.gnd(gnd), .A(_1185_), .Y(_5020_), .vdd(vdd), .B(raddr2_0_bF_buf37_), .C(_5019_), );
  NAND2X1 NAND2X1_965 (.gnd(gnd), .A(regs_24__21_), .Y(_5021_), .vdd(vdd), .B(raddr2_0_bF_buf36_), );
  OAI21X1 OAI21X1_1938 (.gnd(gnd), .A(_3519_), .Y(_5022_), .vdd(vdd), .B(raddr2_0_bF_buf35_), .C(_5021_), );
  MUX2X1 MUX2X1_492 (.gnd(gnd), .A(_5022_), .Y(_5023_), .vdd(vdd), .B(_5020_), .S(raddr2_1_bF_buf1_), );
  MUX2X1 MUX2X1_493 (.gnd(gnd), .A(_5023_), .Y(_5024_), .vdd(vdd), .B(_5018_), .S(raddr2_2_bF_buf9_), );
  MUX2X1 MUX2X1_494 (.gnd(gnd), .A(_5024_), .Y(_5025_), .vdd(vdd), .B(_5015_), .S(_4033__bF_buf3), );
  NAND2X1 NAND2X1_966 (.gnd(gnd), .A(regs_6__21_), .Y(_5026_), .vdd(vdd), .B(raddr2_0_bF_buf34_), );
  OAI21X1 OAI21X1_1939 (.gnd(gnd), .A(_2143_), .Y(_5027_), .vdd(vdd), .B(raddr2_0_bF_buf33_), .C(_5026_), );
  NAND2X1 NAND2X1_967 (.gnd(gnd), .A(regs_4__21_), .Y(_5028_), .vdd(vdd), .B(raddr2_0_bF_buf32_), );
  OAI21X1 OAI21X1_1940 (.gnd(gnd), .A(_3474_), .Y(_5029_), .vdd(vdd), .B(raddr2_0_bF_buf31_), .C(_5028_), );
  MUX2X1 MUX2X1_495 (.gnd(gnd), .A(_5029_), .Y(_5030_), .vdd(vdd), .B(_5027_), .S(raddr2_1_bF_buf0_), );
  NAND2X1 NAND2X1_968 (.gnd(gnd), .A(regs_2__21_), .Y(_5031_), .vdd(vdd), .B(raddr2_0_bF_buf30_), );
  OAI21X1 OAI21X1_1941 (.gnd(gnd), .A(_3483_), .Y(_5032_), .vdd(vdd), .B(raddr2_0_bF_buf29_), .C(_5031_), );
  NAND2X1 NAND2X1_969 (.gnd(gnd), .A(regs_0__21_), .Y(_5033_), .vdd(vdd), .B(raddr2_0_bF_buf28_), );
  OAI21X1 OAI21X1_1942 (.gnd(gnd), .A(_3480_), .Y(_5034_), .vdd(vdd), .B(raddr2_0_bF_buf27_), .C(_5033_), );
  MUX2X1 MUX2X1_496 (.gnd(gnd), .A(_5034_), .Y(_5035_), .vdd(vdd), .B(_5032_), .S(raddr2_1_bF_buf14_bF_buf0_), );
  MUX2X1 MUX2X1_497 (.gnd(gnd), .A(_5035_), .Y(_5036_), .vdd(vdd), .B(_5030_), .S(raddr2_2_bF_buf8_), );
  NAND2X1 NAND2X1_970 (.gnd(gnd), .A(regs_14__21_), .Y(_5037_), .vdd(vdd), .B(raddr2_0_bF_buf26_), );
  OAI21X1 OAI21X1_1943 (.gnd(gnd), .A(_1747_), .Y(_5038_), .vdd(vdd), .B(raddr2_0_bF_buf25_), .C(_5037_), );
  NAND2X1 NAND2X1_971 (.gnd(gnd), .A(regs_12__21_), .Y(_5039_), .vdd(vdd), .B(raddr2_0_bF_buf24_), );
  OAI21X1 OAI21X1_1944 (.gnd(gnd), .A(_1845_), .Y(_5040_), .vdd(vdd), .B(raddr2_0_bF_buf23_), .C(_5039_), );
  MUX2X1 MUX2X1_498 (.gnd(gnd), .A(_5040_), .Y(_5041_), .vdd(vdd), .B(_5038_), .S(raddr2_1_bF_buf13_bF_buf0_), );
  NAND2X1 NAND2X1_972 (.gnd(gnd), .A(regs_10__21_), .Y(_5042_), .vdd(vdd), .B(raddr2_0_bF_buf22_), );
  OAI21X1 OAI21X1_1945 (.gnd(gnd), .A(_1944_), .Y(_5043_), .vdd(vdd), .B(raddr2_0_bF_buf21_), .C(_5042_), );
  NAND2X1 NAND2X1_973 (.gnd(gnd), .A(regs_8__21_), .Y(_5044_), .vdd(vdd), .B(raddr2_0_bF_buf20_), );
  OAI21X1 OAI21X1_1946 (.gnd(gnd), .A(_2042_), .Y(_5045_), .vdd(vdd), .B(raddr2_0_bF_buf19_), .C(_5044_), );
  MUX2X1 MUX2X1_499 (.gnd(gnd), .A(_5045_), .Y(_5046_), .vdd(vdd), .B(_5043_), .S(raddr2_1_bF_buf12_bF_buf0_), );
  MUX2X1 MUX2X1_500 (.gnd(gnd), .A(_5046_), .Y(_5047_), .vdd(vdd), .B(_5041_), .S(raddr2_2_bF_buf7_), );
  MUX2X1 MUX2X1_501 (.gnd(gnd), .A(_5047_), .Y(_5048_), .vdd(vdd), .B(_5036_), .S(_4033__bF_buf2), );
  MUX2X1 MUX2X1_502 (.gnd(gnd), .A(_5048_), .Y(_5512__21_), .vdd(vdd), .B(_5025_), .S(raddr2_4_bF_buf3_), );
  NAND2X1 NAND2X1_974 (.gnd(gnd), .A(regs_22__22_), .Y(_5049_), .vdd(vdd), .B(raddr2_0_bF_buf18_), );
  OAI21X1 OAI21X1_1947 (.gnd(gnd), .A(_1354_), .Y(_5050_), .vdd(vdd), .B(raddr2_0_bF_buf17_), .C(_5049_), );
  NAND2X1 NAND2X1_975 (.gnd(gnd), .A(regs_20__22_), .Y(_5051_), .vdd(vdd), .B(raddr2_0_bF_buf16_), );
  OAI21X1 OAI21X1_1948 (.gnd(gnd), .A(_1452_), .Y(_5052_), .vdd(vdd), .B(raddr2_0_bF_buf15_), .C(_5051_), );
  MUX2X1 MUX2X1_503 (.gnd(gnd), .A(_5052_), .Y(_5053_), .vdd(vdd), .B(_5050_), .S(raddr2_1_bF_buf11_), );
  NAND2X1 NAND2X1_976 (.gnd(gnd), .A(_4036__bF_buf8), .Y(_5054_), .vdd(vdd), .B(_5053_), );
  NAND2X1 NAND2X1_977 (.gnd(gnd), .A(regs_18__22_), .Y(_5055_), .vdd(vdd), .B(raddr2_0_bF_buf14_), );
  OAI21X1 OAI21X1_1949 (.gnd(gnd), .A(_1551_), .Y(_5056_), .vdd(vdd), .B(raddr2_0_bF_buf13_), .C(_5055_), );
  NAND2X1 NAND2X1_978 (.gnd(gnd), .A(regs_16__22_), .Y(_5057_), .vdd(vdd), .B(raddr2_0_bF_buf12_), );
  OAI21X1 OAI21X1_1950 (.gnd(gnd), .A(_1649_), .Y(_5058_), .vdd(vdd), .B(raddr2_0_bF_buf11_), .C(_5057_), );
  MUX2X1 MUX2X1_504 (.gnd(gnd), .A(_5058_), .Y(_5059_), .vdd(vdd), .B(_5056_), .S(raddr2_1_bF_buf10_), );
  AOI21X1 AOI21X1_328 (.gnd(gnd), .A(raddr2_2_bF_buf6_), .Y(_5060_), .vdd(vdd), .B(_5059_), .C(_4033__bF_buf1), );
  OAI21X1 OAI21X1_1951 (.gnd(gnd), .A(_1187_), .Y(_5061_), .vdd(vdd), .B(raddr2_0_bF_buf10_), .C(raddr2_2_bF_buf5_), );
  AOI21X1 AOI21X1_329 (.gnd(gnd), .A(regs_26__22_), .Y(_5062_), .vdd(vdd), .B(raddr2_0_bF_buf9_), .C(_5061_), );
  OAI21X1 OAI21X1_1952 (.gnd(gnd), .A(regs_30__22_), .Y(_5063_), .vdd(vdd), .B(raddr2_2_bF_buf4_), .C(_4038__bF_buf1), );
  OAI21X1 OAI21X1_1953 (.gnd(gnd), .A(_3543_), .Y(_5064_), .vdd(vdd), .B(raddr2_0_bF_buf8_), .C(raddr2_2_bF_buf3_), );
  AOI21X1 AOI21X1_330 (.gnd(gnd), .A(regs_24__22_), .Y(_5065_), .vdd(vdd), .B(raddr2_0_bF_buf7_), .C(_5064_), );
  NOR2X1 NOR2X1_230 (.gnd(gnd), .A(raddr2_0_bF_buf6_), .Y(_5066_), .vdd(vdd), .B(_3537_), );
  NAND2X1 NAND2X1_979 (.gnd(gnd), .A(regs_28__22_), .Y(_5067_), .vdd(vdd), .B(raddr2_0_bF_buf5_), );
  NAND2X1 NAND2X1_980 (.gnd(gnd), .A(_4036__bF_buf7), .Y(_5068_), .vdd(vdd), .B(_5067_), );
  OAI21X1 OAI21X1_1954 (.gnd(gnd), .A(_5068_), .Y(_5069_), .vdd(vdd), .B(_5066_), .C(raddr2_1_bF_buf9_), );
  OAI22X1 OAI22X1_89 (.gnd(gnd), .A(_5062_), .Y(_5070_), .vdd(vdd), .B(_5063_), .C(_5069_), .D(_5065_), );
  AOI22X1 AOI22X1_23 (.gnd(gnd), .A(_5070_), .Y(_5071_), .vdd(vdd), .B(_4033__bF_buf0), .C(_5054_), .D(_5060_), );
  OAI21X1 OAI21X1_1955 (.gnd(gnd), .A(_3551_), .Y(_5072_), .vdd(vdd), .B(raddr2_0_bF_buf4_), .C(raddr2_1_bF_buf8_), );
  AOI21X1 AOI21X1_331 (.gnd(gnd), .A(regs_4__22_), .Y(_5073_), .vdd(vdd), .B(raddr2_0_bF_buf3_), .C(_5072_), );
  AND2X2 AND2X2_68 (.gnd(gnd), .A(regs_6__22_), .Y(_5074_), .vdd(vdd), .B(raddr2_0_bF_buf2_), );
  OAI21X1 OAI21X1_1956 (.gnd(gnd), .A(_2145_), .Y(_5075_), .vdd(vdd), .B(raddr2_0_bF_buf1_), .C(_4038__bF_buf0), );
  OAI21X1 OAI21X1_1957 (.gnd(gnd), .A(_5075_), .Y(_5076_), .vdd(vdd), .B(_5074_), .C(_4036__bF_buf6), );
  OAI21X1 OAI21X1_1958 (.gnd(gnd), .A(_3558_), .Y(_5077_), .vdd(vdd), .B(raddr2_0_bF_buf0_), .C(raddr2_1_bF_buf7_), );
  AOI21X1 AOI21X1_332 (.gnd(gnd), .A(regs_0__22_), .Y(_5078_), .vdd(vdd), .B(raddr2_0_bF_buf96_), .C(_5077_), );
  NOR2X1 NOR2X1_231 (.gnd(gnd), .A(raddr2_0_bF_buf95_), .Y(_5079_), .vdd(vdd), .B(_3555_), );
  NAND2X1 NAND2X1_981 (.gnd(gnd), .A(regs_2__22_), .Y(_5080_), .vdd(vdd), .B(raddr2_0_bF_buf94_), );
  NAND2X1 NAND2X1_982 (.gnd(gnd), .A(_4038__bF_buf8), .Y(_5081_), .vdd(vdd), .B(_5080_), );
  OAI21X1 OAI21X1_1959 (.gnd(gnd), .A(_5081_), .Y(_5082_), .vdd(vdd), .B(_5079_), .C(raddr2_2_bF_buf2_), );
  OAI22X1 OAI22X1_90 (.gnd(gnd), .A(_5078_), .Y(_5083_), .vdd(vdd), .B(_5082_), .C(_5076_), .D(_5073_), );
  NAND2X1 NAND2X1_983 (.gnd(gnd), .A(regs_10__22_), .Y(_5084_), .vdd(vdd), .B(raddr2_0_bF_buf93_), );
  OAI21X1 OAI21X1_1960 (.gnd(gnd), .A(_1946_), .Y(_5085_), .vdd(vdd), .B(raddr2_0_bF_buf92_), .C(_5084_), );
  NAND2X1 NAND2X1_984 (.gnd(gnd), .A(regs_8__22_), .Y(_5086_), .vdd(vdd), .B(raddr2_0_bF_buf91_), );
  OAI21X1 OAI21X1_1961 (.gnd(gnd), .A(_2044_), .Y(_5087_), .vdd(vdd), .B(raddr2_0_bF_buf90_), .C(_5086_), );
  MUX2X1 MUX2X1_505 (.gnd(gnd), .A(_5087_), .Y(_5088_), .vdd(vdd), .B(_5085_), .S(raddr2_1_bF_buf6_), );
  NAND2X1 NAND2X1_985 (.gnd(gnd), .A(regs_14__22_), .Y(_5089_), .vdd(vdd), .B(raddr2_0_bF_buf89_), );
  OAI21X1 OAI21X1_1962 (.gnd(gnd), .A(_1749_), .Y(_5090_), .vdd(vdd), .B(raddr2_0_bF_buf88_), .C(_5089_), );
  NAND2X1 NAND2X1_986 (.gnd(gnd), .A(regs_12__22_), .Y(_5091_), .vdd(vdd), .B(raddr2_0_bF_buf87_), );
  OAI21X1 OAI21X1_1963 (.gnd(gnd), .A(_1847_), .Y(_5092_), .vdd(vdd), .B(raddr2_0_bF_buf86_), .C(_5091_), );
  MUX2X1 MUX2X1_506 (.gnd(gnd), .A(_5092_), .Y(_5093_), .vdd(vdd), .B(_5090_), .S(raddr2_1_bF_buf5_), );
  MUX2X1 MUX2X1_507 (.gnd(gnd), .A(_5093_), .Y(_5094_), .vdd(vdd), .B(_5088_), .S(_4036__bF_buf5), );
  MUX2X1 MUX2X1_508 (.gnd(gnd), .A(_5094_), .Y(_5095_), .vdd(vdd), .B(_5083_), .S(_4033__bF_buf7), );
  MUX2X1 MUX2X1_509 (.gnd(gnd), .A(_5095_), .Y(_5512__22_), .vdd(vdd), .B(_5071_), .S(raddr2_4_bF_buf2_), );
  OAI21X1 OAI21X1_1964 (.gnd(gnd), .A(_1454_), .Y(_5096_), .vdd(vdd), .B(raddr2_0_bF_buf85_), .C(raddr2_1_bF_buf4_), );
  AOI21X1 AOI21X1_333 (.gnd(gnd), .A(regs_20__23_), .Y(_5097_), .vdd(vdd), .B(raddr2_0_bF_buf84_), .C(_5096_), );
  AND2X2 AND2X2_69 (.gnd(gnd), .A(regs_22__23_), .Y(_5098_), .vdd(vdd), .B(raddr2_0_bF_buf83_), );
  OAI21X1 OAI21X1_1965 (.gnd(gnd), .A(_1356_), .Y(_5099_), .vdd(vdd), .B(raddr2_0_bF_buf82_), .C(_4038__bF_buf7), );
  OAI21X1 OAI21X1_1966 (.gnd(gnd), .A(_5099_), .Y(_5100_), .vdd(vdd), .B(_5098_), .C(_4036__bF_buf4), );
  OAI21X1 OAI21X1_1967 (.gnd(gnd), .A(_1651_), .Y(_5101_), .vdd(vdd), .B(raddr2_0_bF_buf81_), .C(raddr2_1_bF_buf3_), );
  AOI21X1 AOI21X1_334 (.gnd(gnd), .A(regs_16__23_), .Y(_5102_), .vdd(vdd), .B(raddr2_0_bF_buf80_), .C(_5101_), );
  NOR2X1 NOR2X1_232 (.gnd(gnd), .A(raddr2_0_bF_buf79_), .Y(_5103_), .vdd(vdd), .B(_1553_), );
  NAND2X1 NAND2X1_987 (.gnd(gnd), .A(regs_18__23_), .Y(_5104_), .vdd(vdd), .B(raddr2_0_bF_buf78_), );
  NAND2X1 NAND2X1_988 (.gnd(gnd), .A(_4038__bF_buf6), .Y(_5105_), .vdd(vdd), .B(_5104_), );
  OAI21X1 OAI21X1_1968 (.gnd(gnd), .A(_5105_), .Y(_5106_), .vdd(vdd), .B(_5103_), .C(raddr2_2_bF_buf1_), );
  OAI22X1 OAI22X1_91 (.gnd(gnd), .A(_5102_), .Y(_5107_), .vdd(vdd), .B(_5106_), .C(_5100_), .D(_5097_), );
  NAND2X1 NAND2X1_989 (.gnd(gnd), .A(regs_28__23_), .Y(_5108_), .vdd(vdd), .B(raddr2_0_bF_buf77_), );
  OAI21X1 OAI21X1_1969 (.gnd(gnd), .A(_3587_), .Y(_5109_), .vdd(vdd), .B(raddr2_0_bF_buf76_), .C(_5108_), );
  MUX2X1 MUX2X1_510 (.gnd(gnd), .A(_5109_), .Y(_5110_), .vdd(vdd), .B(regs_30__23_), .S(raddr2_1_bF_buf2_), );
  NAND2X1 NAND2X1_990 (.gnd(gnd), .A(regs_26__23_), .Y(_5111_), .vdd(vdd), .B(raddr2_0_bF_buf75_), );
  OAI21X1 OAI21X1_1970 (.gnd(gnd), .A(_1189_), .Y(_5112_), .vdd(vdd), .B(raddr2_0_bF_buf74_), .C(_5111_), );
  NAND2X1 NAND2X1_991 (.gnd(gnd), .A(regs_24__23_), .Y(_5113_), .vdd(vdd), .B(raddr2_0_bF_buf73_), );
  OAI21X1 OAI21X1_1971 (.gnd(gnd), .A(_3593_), .Y(_5114_), .vdd(vdd), .B(raddr2_0_bF_buf72_), .C(_5113_), );
  MUX2X1 MUX2X1_511 (.gnd(gnd), .A(_5114_), .Y(_5115_), .vdd(vdd), .B(_5112_), .S(raddr2_1_bF_buf1_), );
  MUX2X1 MUX2X1_512 (.gnd(gnd), .A(_5115_), .Y(_5116_), .vdd(vdd), .B(_5110_), .S(raddr2_2_bF_buf0_), );
  MUX2X1 MUX2X1_513 (.gnd(gnd), .A(_5116_), .Y(_5117_), .vdd(vdd), .B(_5107_), .S(_4033__bF_buf6), );
  NAND2X1 NAND2X1_992 (.gnd(gnd), .A(regs_6__23_), .Y(_5118_), .vdd(vdd), .B(raddr2_0_bF_buf71_), );
  OAI21X1 OAI21X1_1972 (.gnd(gnd), .A(_2147_), .Y(_5119_), .vdd(vdd), .B(raddr2_0_bF_buf70_), .C(_5118_), );
  NAND2X1 NAND2X1_993 (.gnd(gnd), .A(regs_4__23_), .Y(_5120_), .vdd(vdd), .B(raddr2_0_bF_buf69_), );
  OAI21X1 OAI21X1_1973 (.gnd(gnd), .A(_3601_), .Y(_5121_), .vdd(vdd), .B(raddr2_0_bF_buf68_), .C(_5120_), );
  MUX2X1 MUX2X1_514 (.gnd(gnd), .A(_5121_), .Y(_5122_), .vdd(vdd), .B(_5119_), .S(raddr2_1_bF_buf0_), );
  NAND2X1 NAND2X1_994 (.gnd(gnd), .A(regs_2__23_), .Y(_5123_), .vdd(vdd), .B(raddr2_0_bF_buf67_), );
  OAI21X1 OAI21X1_1974 (.gnd(gnd), .A(_3605_), .Y(_5124_), .vdd(vdd), .B(raddr2_0_bF_buf66_), .C(_5123_), );
  NAND2X1 NAND2X1_995 (.gnd(gnd), .A(regs_0__23_), .Y(_5125_), .vdd(vdd), .B(raddr2_0_bF_buf65_), );
  OAI21X1 OAI21X1_1975 (.gnd(gnd), .A(_3608_), .Y(_5126_), .vdd(vdd), .B(raddr2_0_bF_buf64_), .C(_5125_), );
  MUX2X1 MUX2X1_515 (.gnd(gnd), .A(_5126_), .Y(_5127_), .vdd(vdd), .B(_5124_), .S(raddr2_1_bF_buf14_bF_buf3_), );
  MUX2X1 MUX2X1_516 (.gnd(gnd), .A(_5127_), .Y(_5128_), .vdd(vdd), .B(_5122_), .S(raddr2_2_bF_buf10_), );
  NAND2X1 NAND2X1_996 (.gnd(gnd), .A(regs_10__23_), .Y(_5129_), .vdd(vdd), .B(raddr2_0_bF_buf63_), );
  OAI21X1 OAI21X1_1976 (.gnd(gnd), .A(_1948_), .Y(_5130_), .vdd(vdd), .B(raddr2_0_bF_buf62_), .C(_5129_), );
  NAND2X1 NAND2X1_997 (.gnd(gnd), .A(regs_8__23_), .Y(_5131_), .vdd(vdd), .B(raddr2_0_bF_buf61_), );
  OAI21X1 OAI21X1_1977 (.gnd(gnd), .A(_2046_), .Y(_5132_), .vdd(vdd), .B(raddr2_0_bF_buf60_), .C(_5131_), );
  MUX2X1 MUX2X1_517 (.gnd(gnd), .A(_5132_), .Y(_5133_), .vdd(vdd), .B(_5130_), .S(raddr2_1_bF_buf13_bF_buf3_), );
  NAND2X1 NAND2X1_998 (.gnd(gnd), .A(regs_14__23_), .Y(_5134_), .vdd(vdd), .B(raddr2_0_bF_buf59_), );
  OAI21X1 OAI21X1_1978 (.gnd(gnd), .A(_1751_), .Y(_5135_), .vdd(vdd), .B(raddr2_0_bF_buf58_), .C(_5134_), );
  NAND2X1 NAND2X1_999 (.gnd(gnd), .A(regs_12__23_), .Y(_5136_), .vdd(vdd), .B(raddr2_0_bF_buf57_), );
  OAI21X1 OAI21X1_1979 (.gnd(gnd), .A(_1849_), .Y(_5137_), .vdd(vdd), .B(raddr2_0_bF_buf56_), .C(_5136_), );
  MUX2X1 MUX2X1_518 (.gnd(gnd), .A(_5137_), .Y(_5138_), .vdd(vdd), .B(_5135_), .S(raddr2_1_bF_buf12_bF_buf3_), );
  MUX2X1 MUX2X1_519 (.gnd(gnd), .A(_5138_), .Y(_5139_), .vdd(vdd), .B(_5133_), .S(_4036__bF_buf3), );
  MUX2X1 MUX2X1_520 (.gnd(gnd), .A(_5139_), .Y(_5140_), .vdd(vdd), .B(_5128_), .S(_4033__bF_buf5), );
  MUX2X1 MUX2X1_521 (.gnd(gnd), .A(_5140_), .Y(_5512__23_), .vdd(vdd), .B(_5117_), .S(raddr2_4_bF_buf1_), );
  NAND2X1 NAND2X1_1000 (.gnd(gnd), .A(regs_22__24_), .Y(_5141_), .vdd(vdd), .B(raddr2_0_bF_buf55_), );
  OAI21X1 OAI21X1_1980 (.gnd(gnd), .A(_1358_), .Y(_5142_), .vdd(vdd), .B(raddr2_0_bF_buf54_), .C(_5141_), );
  NAND2X1 NAND2X1_1001 (.gnd(gnd), .A(regs_20__24_), .Y(_5143_), .vdd(vdd), .B(raddr2_0_bF_buf53_), );
  OAI21X1 OAI21X1_1981 (.gnd(gnd), .A(_1456_), .Y(_5144_), .vdd(vdd), .B(raddr2_0_bF_buf52_), .C(_5143_), );
  MUX2X1 MUX2X1_522 (.gnd(gnd), .A(_5144_), .Y(_5145_), .vdd(vdd), .B(_5142_), .S(raddr2_1_bF_buf11_), );
  NAND2X1 NAND2X1_1002 (.gnd(gnd), .A(_4036__bF_buf2), .Y(_5146_), .vdd(vdd), .B(_5145_), );
  NAND2X1 NAND2X1_1003 (.gnd(gnd), .A(regs_18__24_), .Y(_5147_), .vdd(vdd), .B(raddr2_0_bF_buf51_), );
  OAI21X1 OAI21X1_1982 (.gnd(gnd), .A(_1555_), .Y(_5148_), .vdd(vdd), .B(raddr2_0_bF_buf50_), .C(_5147_), );
  NAND2X1 NAND2X1_1004 (.gnd(gnd), .A(regs_16__24_), .Y(_5149_), .vdd(vdd), .B(raddr2_0_bF_buf49_), );
  OAI21X1 OAI21X1_1983 (.gnd(gnd), .A(_1653_), .Y(_5150_), .vdd(vdd), .B(raddr2_0_bF_buf48_), .C(_5149_), );
  MUX2X1 MUX2X1_523 (.gnd(gnd), .A(_5150_), .Y(_5151_), .vdd(vdd), .B(_5148_), .S(raddr2_1_bF_buf10_), );
  AOI21X1 AOI21X1_335 (.gnd(gnd), .A(raddr2_2_bF_buf9_), .Y(_5152_), .vdd(vdd), .B(_5151_), .C(_4033__bF_buf4), );
  OAI21X1 OAI21X1_1984 (.gnd(gnd), .A(_1191_), .Y(_5153_), .vdd(vdd), .B(raddr2_0_bF_buf47_), .C(raddr2_2_bF_buf8_), );
  AOI21X1 AOI21X1_336 (.gnd(gnd), .A(regs_26__24_), .Y(_5154_), .vdd(vdd), .B(raddr2_0_bF_buf46_), .C(_5153_), );
  OAI21X1 OAI21X1_1985 (.gnd(gnd), .A(regs_30__24_), .Y(_5155_), .vdd(vdd), .B(raddr2_2_bF_buf7_), .C(_4038__bF_buf5), );
  OAI21X1 OAI21X1_1986 (.gnd(gnd), .A(_3643_), .Y(_5156_), .vdd(vdd), .B(raddr2_0_bF_buf45_), .C(raddr2_2_bF_buf6_), );
  AOI21X1 AOI21X1_337 (.gnd(gnd), .A(regs_24__24_), .Y(_5157_), .vdd(vdd), .B(raddr2_0_bF_buf44_), .C(_5156_), );
  NOR2X1 NOR2X1_233 (.gnd(gnd), .A(raddr2_0_bF_buf43_), .Y(_5158_), .vdd(vdd), .B(_3637_), );
  NAND2X1 NAND2X1_1005 (.gnd(gnd), .A(regs_28__24_), .Y(_5159_), .vdd(vdd), .B(raddr2_0_bF_buf42_), );
  NAND2X1 NAND2X1_1006 (.gnd(gnd), .A(_4036__bF_buf1), .Y(_5160_), .vdd(vdd), .B(_5159_), );
  OAI21X1 OAI21X1_1987 (.gnd(gnd), .A(_5160_), .Y(_5161_), .vdd(vdd), .B(_5158_), .C(raddr2_1_bF_buf9_), );
  OAI22X1 OAI22X1_92 (.gnd(gnd), .A(_5154_), .Y(_5162_), .vdd(vdd), .B(_5155_), .C(_5161_), .D(_5157_), );
  AOI22X1 AOI22X1_24 (.gnd(gnd), .A(_5162_), .Y(_5163_), .vdd(vdd), .B(_4033__bF_buf3), .C(_5146_), .D(_5152_), );
  OAI21X1 OAI21X1_1988 (.gnd(gnd), .A(_3651_), .Y(_5164_), .vdd(vdd), .B(raddr2_0_bF_buf41_), .C(raddr2_1_bF_buf8_), );
  AOI21X1 AOI21X1_338 (.gnd(gnd), .A(regs_4__24_), .Y(_5165_), .vdd(vdd), .B(raddr2_0_bF_buf40_), .C(_5164_), );
  AND2X2 AND2X2_70 (.gnd(gnd), .A(regs_6__24_), .Y(_5166_), .vdd(vdd), .B(raddr2_0_bF_buf39_), );
  OAI21X1 OAI21X1_1989 (.gnd(gnd), .A(_2149_), .Y(_5167_), .vdd(vdd), .B(raddr2_0_bF_buf38_), .C(_4038__bF_buf4), );
  OAI21X1 OAI21X1_1990 (.gnd(gnd), .A(_5167_), .Y(_5168_), .vdd(vdd), .B(_5166_), .C(_4036__bF_buf0), );
  OAI21X1 OAI21X1_1991 (.gnd(gnd), .A(_3658_), .Y(_5169_), .vdd(vdd), .B(raddr2_0_bF_buf37_), .C(raddr2_1_bF_buf7_), );
  AOI21X1 AOI21X1_339 (.gnd(gnd), .A(regs_0__24_), .Y(_5170_), .vdd(vdd), .B(raddr2_0_bF_buf36_), .C(_5169_), );
  NOR2X1 NOR2X1_234 (.gnd(gnd), .A(raddr2_0_bF_buf35_), .Y(_5171_), .vdd(vdd), .B(_3655_), );
  NAND2X1 NAND2X1_1007 (.gnd(gnd), .A(regs_2__24_), .Y(_5172_), .vdd(vdd), .B(raddr2_0_bF_buf34_), );
  NAND2X1 NAND2X1_1008 (.gnd(gnd), .A(_4038__bF_buf3), .Y(_5173_), .vdd(vdd), .B(_5172_), );
  OAI21X1 OAI21X1_1992 (.gnd(gnd), .A(_5173_), .Y(_5174_), .vdd(vdd), .B(_5171_), .C(raddr2_2_bF_buf5_), );
  OAI22X1 OAI22X1_93 (.gnd(gnd), .A(_5170_), .Y(_5175_), .vdd(vdd), .B(_5174_), .C(_5168_), .D(_5165_), );
  NAND2X1 NAND2X1_1009 (.gnd(gnd), .A(regs_10__24_), .Y(_5176_), .vdd(vdd), .B(raddr2_0_bF_buf33_), );
  OAI21X1 OAI21X1_1993 (.gnd(gnd), .A(_1950_), .Y(_5177_), .vdd(vdd), .B(raddr2_0_bF_buf32_), .C(_5176_), );
  NAND2X1 NAND2X1_1010 (.gnd(gnd), .A(regs_8__24_), .Y(_5178_), .vdd(vdd), .B(raddr2_0_bF_buf31_), );
  OAI21X1 OAI21X1_1994 (.gnd(gnd), .A(_2048_), .Y(_5179_), .vdd(vdd), .B(raddr2_0_bF_buf30_), .C(_5178_), );
  MUX2X1 MUX2X1_524 (.gnd(gnd), .A(_5179_), .Y(_5180_), .vdd(vdd), .B(_5177_), .S(raddr2_1_bF_buf6_), );
  NAND2X1 NAND2X1_1011 (.gnd(gnd), .A(regs_14__24_), .Y(_5181_), .vdd(vdd), .B(raddr2_0_bF_buf29_), );
  OAI21X1 OAI21X1_1995 (.gnd(gnd), .A(_1753_), .Y(_5182_), .vdd(vdd), .B(raddr2_0_bF_buf28_), .C(_5181_), );
  NAND2X1 NAND2X1_1012 (.gnd(gnd), .A(regs_12__24_), .Y(_5183_), .vdd(vdd), .B(raddr2_0_bF_buf27_), );
  OAI21X1 OAI21X1_1996 (.gnd(gnd), .A(_1851_), .Y(_5184_), .vdd(vdd), .B(raddr2_0_bF_buf26_), .C(_5183_), );
  MUX2X1 MUX2X1_525 (.gnd(gnd), .A(_5184_), .Y(_5185_), .vdd(vdd), .B(_5182_), .S(raddr2_1_bF_buf5_), );
  MUX2X1 MUX2X1_526 (.gnd(gnd), .A(_5185_), .Y(_5186_), .vdd(vdd), .B(_5180_), .S(_4036__bF_buf8), );
  MUX2X1 MUX2X1_527 (.gnd(gnd), .A(_5186_), .Y(_5187_), .vdd(vdd), .B(_5175_), .S(_4033__bF_buf2), );
  MUX2X1 MUX2X1_528 (.gnd(gnd), .A(_5187_), .Y(_5512__24_), .vdd(vdd), .B(_5163_), .S(raddr2_4_bF_buf0_), );
  NAND2X1 NAND2X1_1013 (.gnd(gnd), .A(regs_22__25_), .Y(_5188_), .vdd(vdd), .B(raddr2_0_bF_buf25_), );
  OAI21X1 OAI21X1_1997 (.gnd(gnd), .A(_1360_), .Y(_5189_), .vdd(vdd), .B(raddr2_0_bF_buf24_), .C(_5188_), );
  NAND2X1 NAND2X1_1014 (.gnd(gnd), .A(regs_20__25_), .Y(_5190_), .vdd(vdd), .B(raddr2_0_bF_buf23_), );
  OAI21X1 OAI21X1_1998 (.gnd(gnd), .A(_1458_), .Y(_5191_), .vdd(vdd), .B(raddr2_0_bF_buf22_), .C(_5190_), );
  MUX2X1 MUX2X1_529 (.gnd(gnd), .A(_5191_), .Y(_5192_), .vdd(vdd), .B(_5189_), .S(raddr2_1_bF_buf4_), );
  NAND2X1 NAND2X1_1015 (.gnd(gnd), .A(_4036__bF_buf7), .Y(_5193_), .vdd(vdd), .B(_5192_), );
  NAND2X1 NAND2X1_1016 (.gnd(gnd), .A(regs_18__25_), .Y(_5194_), .vdd(vdd), .B(raddr2_0_bF_buf21_), );
  OAI21X1 OAI21X1_1999 (.gnd(gnd), .A(_1557_), .Y(_5195_), .vdd(vdd), .B(raddr2_0_bF_buf20_), .C(_5194_), );
  NAND2X1 NAND2X1_1017 (.gnd(gnd), .A(regs_16__25_), .Y(_5196_), .vdd(vdd), .B(raddr2_0_bF_buf19_), );
  OAI21X1 OAI21X1_2000 (.gnd(gnd), .A(_1655_), .Y(_5197_), .vdd(vdd), .B(raddr2_0_bF_buf18_), .C(_5196_), );
  MUX2X1 MUX2X1_530 (.gnd(gnd), .A(_5197_), .Y(_5198_), .vdd(vdd), .B(_5195_), .S(raddr2_1_bF_buf3_), );
  AOI21X1 AOI21X1_340 (.gnd(gnd), .A(raddr2_2_bF_buf4_), .Y(_5199_), .vdd(vdd), .B(_5198_), .C(_4033__bF_buf1), );
  OAI21X1 OAI21X1_2001 (.gnd(gnd), .A(_1193_), .Y(_5200_), .vdd(vdd), .B(raddr2_0_bF_buf17_), .C(raddr2_2_bF_buf3_), );
  AOI21X1 AOI21X1_341 (.gnd(gnd), .A(regs_26__25_), .Y(_5201_), .vdd(vdd), .B(raddr2_0_bF_buf16_), .C(_5200_), );
  OAI21X1 OAI21X1_2002 (.gnd(gnd), .A(regs_30__25_), .Y(_5202_), .vdd(vdd), .B(raddr2_2_bF_buf2_), .C(_4038__bF_buf2), );
  OAI21X1 OAI21X1_2003 (.gnd(gnd), .A(_3720_), .Y(_5203_), .vdd(vdd), .B(raddr2_0_bF_buf15_), .C(raddr2_2_bF_buf1_), );
  AOI21X1 AOI21X1_342 (.gnd(gnd), .A(regs_24__25_), .Y(_5204_), .vdd(vdd), .B(raddr2_0_bF_buf14_), .C(_5203_), );
  NOR2X1 NOR2X1_235 (.gnd(gnd), .A(raddr2_0_bF_buf13_), .Y(_5205_), .vdd(vdd), .B(_3714_), );
  NAND2X1 NAND2X1_1018 (.gnd(gnd), .A(regs_28__25_), .Y(_5206_), .vdd(vdd), .B(raddr2_0_bF_buf12_), );
  NAND2X1 NAND2X1_1019 (.gnd(gnd), .A(_4036__bF_buf6), .Y(_5207_), .vdd(vdd), .B(_5206_), );
  OAI21X1 OAI21X1_2004 (.gnd(gnd), .A(_5207_), .Y(_5208_), .vdd(vdd), .B(_5205_), .C(raddr2_1_bF_buf2_), );
  OAI22X1 OAI22X1_94 (.gnd(gnd), .A(_5201_), .Y(_5209_), .vdd(vdd), .B(_5202_), .C(_5208_), .D(_5204_), );
  AOI22X1 AOI22X1_25 (.gnd(gnd), .A(_5209_), .Y(_5210_), .vdd(vdd), .B(_4033__bF_buf0), .C(_5193_), .D(_5199_), );
  NAND2X1 NAND2X1_1020 (.gnd(gnd), .A(regs_6__25_), .Y(_5211_), .vdd(vdd), .B(raddr2_0_bF_buf11_), );
  OAI21X1 OAI21X1_2005 (.gnd(gnd), .A(_2151_), .Y(_5212_), .vdd(vdd), .B(raddr2_0_bF_buf10_), .C(_5211_), );
  NAND2X1 NAND2X1_1021 (.gnd(gnd), .A(regs_4__25_), .Y(_5213_), .vdd(vdd), .B(raddr2_0_bF_buf9_), );
  OAI21X1 OAI21X1_2006 (.gnd(gnd), .A(_3675_), .Y(_5214_), .vdd(vdd), .B(raddr2_0_bF_buf8_), .C(_5213_), );
  MUX2X1 MUX2X1_531 (.gnd(gnd), .A(_5214_), .Y(_5215_), .vdd(vdd), .B(_5212_), .S(raddr2_1_bF_buf1_), );
  NAND2X1 NAND2X1_1022 (.gnd(gnd), .A(regs_2__25_), .Y(_5216_), .vdd(vdd), .B(raddr2_0_bF_buf7_), );
  OAI21X1 OAI21X1_2007 (.gnd(gnd), .A(_3684_), .Y(_5217_), .vdd(vdd), .B(raddr2_0_bF_buf6_), .C(_5216_), );
  NAND2X1 NAND2X1_1023 (.gnd(gnd), .A(regs_0__25_), .Y(_5218_), .vdd(vdd), .B(raddr2_0_bF_buf5_), );
  OAI21X1 OAI21X1_2008 (.gnd(gnd), .A(_3681_), .Y(_5219_), .vdd(vdd), .B(raddr2_0_bF_buf4_), .C(_5218_), );
  MUX2X1 MUX2X1_532 (.gnd(gnd), .A(_5219_), .Y(_5220_), .vdd(vdd), .B(_5217_), .S(raddr2_1_bF_buf0_), );
  MUX2X1 MUX2X1_533 (.gnd(gnd), .A(_5220_), .Y(_5221_), .vdd(vdd), .B(_5215_), .S(raddr2_2_bF_buf0_), );
  NAND2X1 NAND2X1_1024 (.gnd(gnd), .A(regs_14__25_), .Y(_5222_), .vdd(vdd), .B(raddr2_0_bF_buf3_), );
  OAI21X1 OAI21X1_2009 (.gnd(gnd), .A(_1755_), .Y(_5223_), .vdd(vdd), .B(raddr2_0_bF_buf2_), .C(_5222_), );
  NAND2X1 NAND2X1_1025 (.gnd(gnd), .A(regs_12__25_), .Y(_5224_), .vdd(vdd), .B(raddr2_0_bF_buf1_), );
  OAI21X1 OAI21X1_2010 (.gnd(gnd), .A(_1853_), .Y(_5225_), .vdd(vdd), .B(raddr2_0_bF_buf0_), .C(_5224_), );
  MUX2X1 MUX2X1_534 (.gnd(gnd), .A(_5225_), .Y(_5226_), .vdd(vdd), .B(_5223_), .S(raddr2_1_bF_buf14_bF_buf2_), );
  NAND2X1 NAND2X1_1026 (.gnd(gnd), .A(regs_10__25_), .Y(_5227_), .vdd(vdd), .B(raddr2_0_bF_buf96_), );
  OAI21X1 OAI21X1_2011 (.gnd(gnd), .A(_1952_), .Y(_5228_), .vdd(vdd), .B(raddr2_0_bF_buf95_), .C(_5227_), );
  NAND2X1 NAND2X1_1027 (.gnd(gnd), .A(regs_8__25_), .Y(_5229_), .vdd(vdd), .B(raddr2_0_bF_buf94_), );
  OAI21X1 OAI21X1_2012 (.gnd(gnd), .A(_2050_), .Y(_5230_), .vdd(vdd), .B(raddr2_0_bF_buf93_), .C(_5229_), );
  MUX2X1 MUX2X1_535 (.gnd(gnd), .A(_5230_), .Y(_5231_), .vdd(vdd), .B(_5228_), .S(raddr2_1_bF_buf13_bF_buf2_), );
  MUX2X1 MUX2X1_536 (.gnd(gnd), .A(_5231_), .Y(_5232_), .vdd(vdd), .B(_5226_), .S(raddr2_2_bF_buf10_), );
  MUX2X1 MUX2X1_537 (.gnd(gnd), .A(_5232_), .Y(_5233_), .vdd(vdd), .B(_5221_), .S(_4033__bF_buf7), );
  MUX2X1 MUX2X1_538 (.gnd(gnd), .A(_5233_), .Y(_5512__25_), .vdd(vdd), .B(_5210_), .S(raddr2_4_bF_buf4_), );
  OAI21X1 OAI21X1_2013 (.gnd(gnd), .A(_3726_), .Y(_5234_), .vdd(vdd), .B(raddr2_0_bF_buf92_), .C(raddr2_1_bF_buf12_bF_buf2_), );
  AOI21X1 AOI21X1_343 (.gnd(gnd), .A(regs_4__26_), .Y(_5235_), .vdd(vdd), .B(raddr2_0_bF_buf91_), .C(_5234_), );
  AND2X2 AND2X2_71 (.gnd(gnd), .A(regs_6__26_), .Y(_5236_), .vdd(vdd), .B(raddr2_0_bF_buf90_), );
  OAI21X1 OAI21X1_2014 (.gnd(gnd), .A(_2153_), .Y(_5237_), .vdd(vdd), .B(raddr2_0_bF_buf89_), .C(_4038__bF_buf1), );
  OAI21X1 OAI21X1_2015 (.gnd(gnd), .A(_5237_), .Y(_5238_), .vdd(vdd), .B(_5236_), .C(_4036__bF_buf5), );
  OAI21X1 OAI21X1_2016 (.gnd(gnd), .A(_3732_), .Y(_5239_), .vdd(vdd), .B(raddr2_0_bF_buf88_), .C(raddr2_1_bF_buf11_), );
  AOI21X1 AOI21X1_344 (.gnd(gnd), .A(regs_0__26_), .Y(_5240_), .vdd(vdd), .B(raddr2_0_bF_buf87_), .C(_5239_), );
  NOR2X1 NOR2X1_236 (.gnd(gnd), .A(raddr2_0_bF_buf86_), .Y(_5241_), .vdd(vdd), .B(_3735_), );
  NAND2X1 NAND2X1_1028 (.gnd(gnd), .A(regs_2__26_), .Y(_5242_), .vdd(vdd), .B(raddr2_0_bF_buf85_), );
  NAND2X1 NAND2X1_1029 (.gnd(gnd), .A(_4038__bF_buf0), .Y(_5243_), .vdd(vdd), .B(_5242_), );
  OAI21X1 OAI21X1_2017 (.gnd(gnd), .A(_5243_), .Y(_5244_), .vdd(vdd), .B(_5241_), .C(raddr2_2_bF_buf9_), );
  OAI22X1 OAI22X1_95 (.gnd(gnd), .A(_5240_), .Y(_5245_), .vdd(vdd), .B(_5244_), .C(_5238_), .D(_5235_), );
  NAND2X1 NAND2X1_1030 (.gnd(gnd), .A(regs_10__26_), .Y(_5246_), .vdd(vdd), .B(raddr2_0_bF_buf84_), );
  OAI21X1 OAI21X1_2018 (.gnd(gnd), .A(_1954_), .Y(_5247_), .vdd(vdd), .B(raddr2_0_bF_buf83_), .C(_5246_), );
  NAND2X1 NAND2X1_1031 (.gnd(gnd), .A(regs_8__26_), .Y(_5248_), .vdd(vdd), .B(raddr2_0_bF_buf82_), );
  OAI21X1 OAI21X1_2019 (.gnd(gnd), .A(_2052_), .Y(_5249_), .vdd(vdd), .B(raddr2_0_bF_buf81_), .C(_5248_), );
  MUX2X1 MUX2X1_539 (.gnd(gnd), .A(_5249_), .Y(_5250_), .vdd(vdd), .B(_5247_), .S(raddr2_1_bF_buf10_), );
  NAND2X1 NAND2X1_1032 (.gnd(gnd), .A(regs_14__26_), .Y(_5251_), .vdd(vdd), .B(raddr2_0_bF_buf80_), );
  OAI21X1 OAI21X1_2020 (.gnd(gnd), .A(_1757_), .Y(_5252_), .vdd(vdd), .B(raddr2_0_bF_buf79_), .C(_5251_), );
  NAND2X1 NAND2X1_1033 (.gnd(gnd), .A(regs_12__26_), .Y(_5253_), .vdd(vdd), .B(raddr2_0_bF_buf78_), );
  OAI21X1 OAI21X1_2021 (.gnd(gnd), .A(_1855_), .Y(_5254_), .vdd(vdd), .B(raddr2_0_bF_buf77_), .C(_5253_), );
  MUX2X1 MUX2X1_540 (.gnd(gnd), .A(_5254_), .Y(_5255_), .vdd(vdd), .B(_5252_), .S(raddr2_1_bF_buf9_), );
  MUX2X1 MUX2X1_541 (.gnd(gnd), .A(_5255_), .Y(_5256_), .vdd(vdd), .B(_5250_), .S(_4036__bF_buf4), );
  MUX2X1 MUX2X1_542 (.gnd(gnd), .A(_5256_), .Y(_5257_), .vdd(vdd), .B(_5245_), .S(_4033__bF_buf6), );
  OAI21X1 OAI21X1_2022 (.gnd(gnd), .A(_1657_), .Y(_5258_), .vdd(vdd), .B(raddr2_0_bF_buf76_), .C(raddr2_1_bF_buf8_), );
  AOI21X1 AOI21X1_345 (.gnd(gnd), .A(regs_16__26_), .Y(_5259_), .vdd(vdd), .B(raddr2_0_bF_buf75_), .C(_5258_), );
  NOR2X1 NOR2X1_237 (.gnd(gnd), .A(raddr2_0_bF_buf74_), .Y(_5260_), .vdd(vdd), .B(_1559_), );
  NAND2X1 NAND2X1_1034 (.gnd(gnd), .A(regs_18__26_), .Y(_5261_), .vdd(vdd), .B(raddr2_0_bF_buf73_), );
  NAND2X1 NAND2X1_1035 (.gnd(gnd), .A(_4038__bF_buf8), .Y(_5262_), .vdd(vdd), .B(_5261_), );
  OAI21X1 OAI21X1_2023 (.gnd(gnd), .A(_5262_), .Y(_5263_), .vdd(vdd), .B(_5260_), .C(raddr2_2_bF_buf8_), );
  OAI21X1 OAI21X1_2024 (.gnd(gnd), .A(_1460_), .Y(_5264_), .vdd(vdd), .B(raddr2_0_bF_buf72_), .C(raddr2_1_bF_buf7_), );
  AOI21X1 AOI21X1_346 (.gnd(gnd), .A(regs_20__26_), .Y(_5265_), .vdd(vdd), .B(raddr2_0_bF_buf71_), .C(_5264_), );
  AND2X2 AND2X2_72 (.gnd(gnd), .A(regs_22__26_), .Y(_5266_), .vdd(vdd), .B(raddr2_0_bF_buf70_), );
  OAI21X1 OAI21X1_2025 (.gnd(gnd), .A(_1362_), .Y(_5267_), .vdd(vdd), .B(raddr2_0_bF_buf69_), .C(_4038__bF_buf7), );
  OAI21X1 OAI21X1_2026 (.gnd(gnd), .A(_5267_), .Y(_5268_), .vdd(vdd), .B(_5266_), .C(_4036__bF_buf3), );
  OAI22X1 OAI22X1_96 (.gnd(gnd), .A(_5259_), .Y(_5269_), .vdd(vdd), .B(_5263_), .C(_5268_), .D(_5265_), );
  NAND2X1 NAND2X1_1036 (.gnd(gnd), .A(regs_28__26_), .Y(_5270_), .vdd(vdd), .B(raddr2_0_bF_buf68_), );
  OAI21X1 OAI21X1_2027 (.gnd(gnd), .A(_3765_), .Y(_5271_), .vdd(vdd), .B(raddr2_0_bF_buf67_), .C(_5270_), );
  MUX2X1 MUX2X1_543 (.gnd(gnd), .A(_5271_), .Y(_5272_), .vdd(vdd), .B(regs_30__26_), .S(raddr2_1_bF_buf6_), );
  NAND2X1 NAND2X1_1037 (.gnd(gnd), .A(regs_26__26_), .Y(_5273_), .vdd(vdd), .B(raddr2_0_bF_buf66_), );
  OAI21X1 OAI21X1_2028 (.gnd(gnd), .A(_1195_), .Y(_5274_), .vdd(vdd), .B(raddr2_0_bF_buf65_), .C(_5273_), );
  NAND2X1 NAND2X1_1038 (.gnd(gnd), .A(regs_24__26_), .Y(_5275_), .vdd(vdd), .B(raddr2_0_bF_buf64_), );
  OAI21X1 OAI21X1_2029 (.gnd(gnd), .A(_3771_), .Y(_5276_), .vdd(vdd), .B(raddr2_0_bF_buf63_), .C(_5275_), );
  MUX2X1 MUX2X1_544 (.gnd(gnd), .A(_5276_), .Y(_5277_), .vdd(vdd), .B(_5274_), .S(raddr2_1_bF_buf5_), );
  MUX2X1 MUX2X1_545 (.gnd(gnd), .A(_5277_), .Y(_5278_), .vdd(vdd), .B(_5272_), .S(raddr2_2_bF_buf7_), );
  MUX2X1 MUX2X1_546 (.gnd(gnd), .A(_5278_), .Y(_5279_), .vdd(vdd), .B(_5269_), .S(_4033__bF_buf5), );
  MUX2X1 MUX2X1_547 (.gnd(gnd), .A(_5257_), .Y(_5512__26_), .vdd(vdd), .B(_5279_), .S(raddr2_4_bF_buf3_), );
  OAI21X1 OAI21X1_2030 (.gnd(gnd), .A(_1462_), .Y(_5280_), .vdd(vdd), .B(raddr2_0_bF_buf62_), .C(raddr2_1_bF_buf4_), );
  AOI21X1 AOI21X1_347 (.gnd(gnd), .A(regs_20__27_), .Y(_5281_), .vdd(vdd), .B(raddr2_0_bF_buf61_), .C(_5280_), );
  AND2X2 AND2X2_73 (.gnd(gnd), .A(regs_22__27_), .Y(_5282_), .vdd(vdd), .B(raddr2_0_bF_buf60_), );
  OAI21X1 OAI21X1_2031 (.gnd(gnd), .A(_1364_), .Y(_5283_), .vdd(vdd), .B(raddr2_0_bF_buf59_), .C(_4038__bF_buf6), );
  OAI21X1 OAI21X1_2032 (.gnd(gnd), .A(_5283_), .Y(_5284_), .vdd(vdd), .B(_5282_), .C(_4036__bF_buf2), );
  OAI21X1 OAI21X1_2033 (.gnd(gnd), .A(_1659_), .Y(_5285_), .vdd(vdd), .B(raddr2_0_bF_buf58_), .C(raddr2_1_bF_buf3_), );
  AOI21X1 AOI21X1_348 (.gnd(gnd), .A(regs_16__27_), .Y(_5286_), .vdd(vdd), .B(raddr2_0_bF_buf57_), .C(_5285_), );
  NOR2X1 NOR2X1_238 (.gnd(gnd), .A(raddr2_0_bF_buf56_), .Y(_5287_), .vdd(vdd), .B(_1561_), );
  NAND2X1 NAND2X1_1039 (.gnd(gnd), .A(regs_18__27_), .Y(_5288_), .vdd(vdd), .B(raddr2_0_bF_buf55_), );
  NAND2X1 NAND2X1_1040 (.gnd(gnd), .A(_4038__bF_buf5), .Y(_5289_), .vdd(vdd), .B(_5288_), );
  OAI21X1 OAI21X1_2034 (.gnd(gnd), .A(_5289_), .Y(_5290_), .vdd(vdd), .B(_5287_), .C(raddr2_2_bF_buf6_), );
  OAI22X1 OAI22X1_97 (.gnd(gnd), .A(_5286_), .Y(_5291_), .vdd(vdd), .B(_5290_), .C(_5284_), .D(_5281_), );
  NAND2X1 NAND2X1_1041 (.gnd(gnd), .A(regs_28__27_), .Y(_5292_), .vdd(vdd), .B(raddr2_0_bF_buf54_), );
  OAI21X1 OAI21X1_2035 (.gnd(gnd), .A(_3795_), .Y(_5293_), .vdd(vdd), .B(raddr2_0_bF_buf53_), .C(_5292_), );
  MUX2X1 MUX2X1_548 (.gnd(gnd), .A(_5293_), .Y(_5294_), .vdd(vdd), .B(regs_30__27_), .S(raddr2_1_bF_buf2_), );
  NAND2X1 NAND2X1_1042 (.gnd(gnd), .A(regs_26__27_), .Y(_5295_), .vdd(vdd), .B(raddr2_0_bF_buf52_), );
  OAI21X1 OAI21X1_2036 (.gnd(gnd), .A(_1197_), .Y(_5296_), .vdd(vdd), .B(raddr2_0_bF_buf51_), .C(_5295_), );
  NAND2X1 NAND2X1_1043 (.gnd(gnd), .A(regs_24__27_), .Y(_5297_), .vdd(vdd), .B(raddr2_0_bF_buf50_), );
  OAI21X1 OAI21X1_2037 (.gnd(gnd), .A(_3792_), .Y(_5298_), .vdd(vdd), .B(raddr2_0_bF_buf49_), .C(_5297_), );
  MUX2X1 MUX2X1_549 (.gnd(gnd), .A(_5298_), .Y(_5299_), .vdd(vdd), .B(_5296_), .S(raddr2_1_bF_buf1_), );
  MUX2X1 MUX2X1_550 (.gnd(gnd), .A(_5299_), .Y(_5300_), .vdd(vdd), .B(_5294_), .S(raddr2_2_bF_buf5_), );
  MUX2X1 MUX2X1_551 (.gnd(gnd), .A(_5300_), .Y(_5301_), .vdd(vdd), .B(_5291_), .S(_4033__bF_buf4), );
  NAND2X1 NAND2X1_1044 (.gnd(gnd), .A(regs_6__27_), .Y(_5302_), .vdd(vdd), .B(raddr2_0_bF_buf48_), );
  OAI21X1 OAI21X1_2038 (.gnd(gnd), .A(_2155_), .Y(_5303_), .vdd(vdd), .B(raddr2_0_bF_buf47_), .C(_5302_), );
  NAND2X1 NAND2X1_1045 (.gnd(gnd), .A(regs_4__27_), .Y(_5304_), .vdd(vdd), .B(raddr2_0_bF_buf46_), );
  OAI21X1 OAI21X1_2039 (.gnd(gnd), .A(_3804_), .Y(_5305_), .vdd(vdd), .B(raddr2_0_bF_buf45_), .C(_5304_), );
  MUX2X1 MUX2X1_552 (.gnd(gnd), .A(_5305_), .Y(_5306_), .vdd(vdd), .B(_5303_), .S(raddr2_1_bF_buf0_), );
  NAND2X1 NAND2X1_1046 (.gnd(gnd), .A(regs_2__27_), .Y(_5307_), .vdd(vdd), .B(raddr2_0_bF_buf44_), );
  OAI21X1 OAI21X1_2040 (.gnd(gnd), .A(_3808_), .Y(_5308_), .vdd(vdd), .B(raddr2_0_bF_buf43_), .C(_5307_), );
  NAND2X1 NAND2X1_1047 (.gnd(gnd), .A(regs_0__27_), .Y(_5309_), .vdd(vdd), .B(raddr2_0_bF_buf42_), );
  OAI21X1 OAI21X1_2041 (.gnd(gnd), .A(_3811_), .Y(_5310_), .vdd(vdd), .B(raddr2_0_bF_buf41_), .C(_5309_), );
  MUX2X1 MUX2X1_553 (.gnd(gnd), .A(_5310_), .Y(_5311_), .vdd(vdd), .B(_5308_), .S(raddr2_1_bF_buf14_bF_buf1_), );
  MUX2X1 MUX2X1_554 (.gnd(gnd), .A(_5311_), .Y(_5312_), .vdd(vdd), .B(_5306_), .S(raddr2_2_bF_buf4_), );
  NAND2X1 NAND2X1_1048 (.gnd(gnd), .A(regs_10__27_), .Y(_5313_), .vdd(vdd), .B(raddr2_0_bF_buf40_), );
  OAI21X1 OAI21X1_2042 (.gnd(gnd), .A(_1956_), .Y(_5314_), .vdd(vdd), .B(raddr2_0_bF_buf39_), .C(_5313_), );
  NAND2X1 NAND2X1_1049 (.gnd(gnd), .A(regs_8__27_), .Y(_5315_), .vdd(vdd), .B(raddr2_0_bF_buf38_), );
  OAI21X1 OAI21X1_2043 (.gnd(gnd), .A(_2054_), .Y(_5316_), .vdd(vdd), .B(raddr2_0_bF_buf37_), .C(_5315_), );
  MUX2X1 MUX2X1_555 (.gnd(gnd), .A(_5316_), .Y(_5317_), .vdd(vdd), .B(_5314_), .S(raddr2_1_bF_buf13_bF_buf1_), );
  NAND2X1 NAND2X1_1050 (.gnd(gnd), .A(regs_14__27_), .Y(_5318_), .vdd(vdd), .B(raddr2_0_bF_buf36_), );
  OAI21X1 OAI21X1_2044 (.gnd(gnd), .A(_1759_), .Y(_5319_), .vdd(vdd), .B(raddr2_0_bF_buf35_), .C(_5318_), );
  NAND2X1 NAND2X1_1051 (.gnd(gnd), .A(regs_12__27_), .Y(_5320_), .vdd(vdd), .B(raddr2_0_bF_buf34_), );
  OAI21X1 OAI21X1_2045 (.gnd(gnd), .A(_1857_), .Y(_5321_), .vdd(vdd), .B(raddr2_0_bF_buf33_), .C(_5320_), );
  MUX2X1 MUX2X1_556 (.gnd(gnd), .A(_5321_), .Y(_5322_), .vdd(vdd), .B(_5319_), .S(raddr2_1_bF_buf12_bF_buf1_), );
  MUX2X1 MUX2X1_557 (.gnd(gnd), .A(_5322_), .Y(_5323_), .vdd(vdd), .B(_5317_), .S(_4036__bF_buf1), );
  MUX2X1 MUX2X1_558 (.gnd(gnd), .A(_5323_), .Y(_5324_), .vdd(vdd), .B(_5312_), .S(_4033__bF_buf3), );
  MUX2X1 MUX2X1_559 (.gnd(gnd), .A(_5324_), .Y(_5512__27_), .vdd(vdd), .B(_5301_), .S(raddr2_4_bF_buf2_), );
  NAND2X1 NAND2X1_1052 (.gnd(gnd), .A(regs_22__28_), .Y(_5325_), .vdd(vdd), .B(raddr2_0_bF_buf32_), );
  OAI21X1 OAI21X1_2046 (.gnd(gnd), .A(_1366_), .Y(_5326_), .vdd(vdd), .B(raddr2_0_bF_buf31_), .C(_5325_), );
  NAND2X1 NAND2X1_1053 (.gnd(gnd), .A(regs_20__28_), .Y(_5327_), .vdd(vdd), .B(raddr2_0_bF_buf30_), );
  OAI21X1 OAI21X1_2047 (.gnd(gnd), .A(_1464_), .Y(_5328_), .vdd(vdd), .B(raddr2_0_bF_buf29_), .C(_5327_), );
  MUX2X1 MUX2X1_560 (.gnd(gnd), .A(_5328_), .Y(_5329_), .vdd(vdd), .B(_5326_), .S(raddr2_1_bF_buf11_), );
  NAND2X1 NAND2X1_1054 (.gnd(gnd), .A(_4036__bF_buf0), .Y(_5330_), .vdd(vdd), .B(_5329_), );
  NAND2X1 NAND2X1_1055 (.gnd(gnd), .A(regs_18__28_), .Y(_5331_), .vdd(vdd), .B(raddr2_0_bF_buf28_), );
  OAI21X1 OAI21X1_2048 (.gnd(gnd), .A(_1563_), .Y(_5332_), .vdd(vdd), .B(raddr2_0_bF_buf27_), .C(_5331_), );
  NAND2X1 NAND2X1_1056 (.gnd(gnd), .A(regs_16__28_), .Y(_5333_), .vdd(vdd), .B(raddr2_0_bF_buf26_), );
  OAI21X1 OAI21X1_2049 (.gnd(gnd), .A(_1661_), .Y(_5334_), .vdd(vdd), .B(raddr2_0_bF_buf25_), .C(_5333_), );
  MUX2X1 MUX2X1_561 (.gnd(gnd), .A(_5334_), .Y(_5335_), .vdd(vdd), .B(_5332_), .S(raddr2_1_bF_buf10_), );
  AOI21X1 AOI21X1_349 (.gnd(gnd), .A(raddr2_2_bF_buf3_), .Y(_5336_), .vdd(vdd), .B(_5335_), .C(_4033__bF_buf2), );
  OAI21X1 OAI21X1_2050 (.gnd(gnd), .A(_1199_), .Y(_5337_), .vdd(vdd), .B(raddr2_0_bF_buf24_), .C(raddr2_2_bF_buf2_), );
  AOI21X1 AOI21X1_350 (.gnd(gnd), .A(regs_26__28_), .Y(_5338_), .vdd(vdd), .B(raddr2_0_bF_buf23_), .C(_5337_), );
  OAI21X1 OAI21X1_2051 (.gnd(gnd), .A(regs_30__28_), .Y(_5339_), .vdd(vdd), .B(raddr2_2_bF_buf1_), .C(_4038__bF_buf4), );
  OAI21X1 OAI21X1_2052 (.gnd(gnd), .A(_3843_), .Y(_5340_), .vdd(vdd), .B(raddr2_0_bF_buf22_), .C(raddr2_2_bF_buf0_), );
  AOI21X1 AOI21X1_351 (.gnd(gnd), .A(regs_24__28_), .Y(_5341_), .vdd(vdd), .B(raddr2_0_bF_buf21_), .C(_5340_), );
  NOR2X1 NOR2X1_239 (.gnd(gnd), .A(raddr2_0_bF_buf20_), .Y(_5342_), .vdd(vdd), .B(_3846_), );
  NAND2X1 NAND2X1_1057 (.gnd(gnd), .A(regs_28__28_), .Y(_5343_), .vdd(vdd), .B(raddr2_0_bF_buf19_), );
  NAND2X1 NAND2X1_1058 (.gnd(gnd), .A(_4036__bF_buf8), .Y(_5344_), .vdd(vdd), .B(_5343_), );
  OAI21X1 OAI21X1_2053 (.gnd(gnd), .A(_5344_), .Y(_5345_), .vdd(vdd), .B(_5342_), .C(raddr2_1_bF_buf9_), );
  OAI22X1 OAI22X1_98 (.gnd(gnd), .A(_5338_), .Y(_5346_), .vdd(vdd), .B(_5339_), .C(_5345_), .D(_5341_), );
  AOI22X1 AOI22X1_26 (.gnd(gnd), .A(_5346_), .Y(_5347_), .vdd(vdd), .B(_4033__bF_buf1), .C(_5330_), .D(_5336_), );
  OAI21X1 OAI21X1_2054 (.gnd(gnd), .A(_3853_), .Y(_5348_), .vdd(vdd), .B(raddr2_0_bF_buf18_), .C(raddr2_1_bF_buf8_), );
  AOI21X1 AOI21X1_352 (.gnd(gnd), .A(regs_4__28_), .Y(_5349_), .vdd(vdd), .B(raddr2_0_bF_buf17_), .C(_5348_), );
  AND2X2 AND2X2_74 (.gnd(gnd), .A(regs_6__28_), .Y(_5350_), .vdd(vdd), .B(raddr2_0_bF_buf16_), );
  OAI21X1 OAI21X1_2055 (.gnd(gnd), .A(_2157_), .Y(_5351_), .vdd(vdd), .B(raddr2_0_bF_buf15_), .C(_4038__bF_buf3), );
  OAI21X1 OAI21X1_2056 (.gnd(gnd), .A(_5351_), .Y(_5352_), .vdd(vdd), .B(_5350_), .C(_4036__bF_buf7), );
  OAI21X1 OAI21X1_2057 (.gnd(gnd), .A(_3859_), .Y(_5353_), .vdd(vdd), .B(raddr2_0_bF_buf14_), .C(raddr2_1_bF_buf7_), );
  AOI21X1 AOI21X1_353 (.gnd(gnd), .A(regs_0__28_), .Y(_5354_), .vdd(vdd), .B(raddr2_0_bF_buf13_), .C(_5353_), );
  NOR2X1 NOR2X1_240 (.gnd(gnd), .A(raddr2_0_bF_buf12_), .Y(_5355_), .vdd(vdd), .B(_3862_), );
  NAND2X1 NAND2X1_1059 (.gnd(gnd), .A(regs_2__28_), .Y(_5356_), .vdd(vdd), .B(raddr2_0_bF_buf11_), );
  NAND2X1 NAND2X1_1060 (.gnd(gnd), .A(_4038__bF_buf2), .Y(_5357_), .vdd(vdd), .B(_5356_), );
  OAI21X1 OAI21X1_2058 (.gnd(gnd), .A(_5357_), .Y(_5358_), .vdd(vdd), .B(_5355_), .C(raddr2_2_bF_buf10_), );
  OAI22X1 OAI22X1_99 (.gnd(gnd), .A(_5354_), .Y(_5359_), .vdd(vdd), .B(_5358_), .C(_5352_), .D(_5349_), );
  NAND2X1 NAND2X1_1061 (.gnd(gnd), .A(regs_10__28_), .Y(_5360_), .vdd(vdd), .B(raddr2_0_bF_buf10_), );
  OAI21X1 OAI21X1_2059 (.gnd(gnd), .A(_1958_), .Y(_5361_), .vdd(vdd), .B(raddr2_0_bF_buf9_), .C(_5360_), );
  NAND2X1 NAND2X1_1062 (.gnd(gnd), .A(regs_8__28_), .Y(_5362_), .vdd(vdd), .B(raddr2_0_bF_buf8_), );
  OAI21X1 OAI21X1_2060 (.gnd(gnd), .A(_2056_), .Y(_5363_), .vdd(vdd), .B(raddr2_0_bF_buf7_), .C(_5362_), );
  MUX2X1 MUX2X1_562 (.gnd(gnd), .A(_5363_), .Y(_5364_), .vdd(vdd), .B(_5361_), .S(raddr2_1_bF_buf6_), );
  NAND2X1 NAND2X1_1063 (.gnd(gnd), .A(regs_14__28_), .Y(_5365_), .vdd(vdd), .B(raddr2_0_bF_buf6_), );
  OAI21X1 OAI21X1_2061 (.gnd(gnd), .A(_1761_), .Y(_5366_), .vdd(vdd), .B(raddr2_0_bF_buf5_), .C(_5365_), );
  NAND2X1 NAND2X1_1064 (.gnd(gnd), .A(regs_12__28_), .Y(_5367_), .vdd(vdd), .B(raddr2_0_bF_buf4_), );
  OAI21X1 OAI21X1_2062 (.gnd(gnd), .A(_1859_), .Y(_5368_), .vdd(vdd), .B(raddr2_0_bF_buf3_), .C(_5367_), );
  MUX2X1 MUX2X1_563 (.gnd(gnd), .A(_5368_), .Y(_5369_), .vdd(vdd), .B(_5366_), .S(raddr2_1_bF_buf5_), );
  MUX2X1 MUX2X1_564 (.gnd(gnd), .A(_5369_), .Y(_5370_), .vdd(vdd), .B(_5364_), .S(_4036__bF_buf6), );
  MUX2X1 MUX2X1_565 (.gnd(gnd), .A(_5370_), .Y(_5371_), .vdd(vdd), .B(_5359_), .S(_4033__bF_buf0), );
  MUX2X1 MUX2X1_566 (.gnd(gnd), .A(_5371_), .Y(_5512__28_), .vdd(vdd), .B(_5347_), .S(raddr2_4_bF_buf1_), );
  OAI21X1 OAI21X1_2063 (.gnd(gnd), .A(_3905_), .Y(_5372_), .vdd(vdd), .B(raddr2_0_bF_buf2_), .C(raddr2_1_bF_buf4_), );
  AOI21X1 AOI21X1_354 (.gnd(gnd), .A(regs_4__29_), .Y(_5373_), .vdd(vdd), .B(raddr2_0_bF_buf1_), .C(_5372_), );
  AND2X2 AND2X2_75 (.gnd(gnd), .A(regs_6__29_), .Y(_5374_), .vdd(vdd), .B(raddr2_0_bF_buf0_), );
  OAI21X1 OAI21X1_2064 (.gnd(gnd), .A(_2159_), .Y(_5375_), .vdd(vdd), .B(raddr2_0_bF_buf96_), .C(_4038__bF_buf1), );
  OAI21X1 OAI21X1_2065 (.gnd(gnd), .A(_5375_), .Y(_5376_), .vdd(vdd), .B(_5374_), .C(_4036__bF_buf5), );
  OAI21X1 OAI21X1_2066 (.gnd(gnd), .A(_3911_), .Y(_5377_), .vdd(vdd), .B(raddr2_0_bF_buf95_), .C(raddr2_1_bF_buf3_), );
  AOI21X1 AOI21X1_355 (.gnd(gnd), .A(regs_0__29_), .Y(_5378_), .vdd(vdd), .B(raddr2_0_bF_buf94_), .C(_5377_), );
  NOR2X1 NOR2X1_241 (.gnd(gnd), .A(raddr2_0_bF_buf93_), .Y(_5379_), .vdd(vdd), .B(_3914_), );
  NAND2X1 NAND2X1_1065 (.gnd(gnd), .A(regs_2__29_), .Y(_5380_), .vdd(vdd), .B(raddr2_0_bF_buf92_), );
  NAND2X1 NAND2X1_1066 (.gnd(gnd), .A(_4038__bF_buf0), .Y(_5381_), .vdd(vdd), .B(_5380_), );
  OAI21X1 OAI21X1_2067 (.gnd(gnd), .A(_5381_), .Y(_5382_), .vdd(vdd), .B(_5379_), .C(raddr2_2_bF_buf9_), );
  OAI22X1 OAI22X1_100 (.gnd(gnd), .A(_5378_), .Y(_5383_), .vdd(vdd), .B(_5382_), .C(_5376_), .D(_5373_), );
  NAND2X1 NAND2X1_1067 (.gnd(gnd), .A(regs_10__29_), .Y(_5384_), .vdd(vdd), .B(raddr2_0_bF_buf91_), );
  OAI21X1 OAI21X1_2068 (.gnd(gnd), .A(_1960_), .Y(_5385_), .vdd(vdd), .B(raddr2_0_bF_buf90_), .C(_5384_), );
  NAND2X1 NAND2X1_1068 (.gnd(gnd), .A(regs_8__29_), .Y(_5386_), .vdd(vdd), .B(raddr2_0_bF_buf89_), );
  OAI21X1 OAI21X1_2069 (.gnd(gnd), .A(_2058_), .Y(_5387_), .vdd(vdd), .B(raddr2_0_bF_buf88_), .C(_5386_), );
  MUX2X1 MUX2X1_567 (.gnd(gnd), .A(_5387_), .Y(_5388_), .vdd(vdd), .B(_5385_), .S(raddr2_1_bF_buf2_), );
  NAND2X1 NAND2X1_1069 (.gnd(gnd), .A(regs_14__29_), .Y(_5389_), .vdd(vdd), .B(raddr2_0_bF_buf87_), );
  OAI21X1 OAI21X1_2070 (.gnd(gnd), .A(_1763_), .Y(_5390_), .vdd(vdd), .B(raddr2_0_bF_buf86_), .C(_5389_), );
  NAND2X1 NAND2X1_1070 (.gnd(gnd), .A(regs_12__29_), .Y(_5391_), .vdd(vdd), .B(raddr2_0_bF_buf85_), );
  OAI21X1 OAI21X1_2071 (.gnd(gnd), .A(_1861_), .Y(_5392_), .vdd(vdd), .B(raddr2_0_bF_buf84_), .C(_5391_), );
  MUX2X1 MUX2X1_568 (.gnd(gnd), .A(_5392_), .Y(_5393_), .vdd(vdd), .B(_5390_), .S(raddr2_1_bF_buf1_), );
  MUX2X1 MUX2X1_569 (.gnd(gnd), .A(_5393_), .Y(_5394_), .vdd(vdd), .B(_5388_), .S(_4036__bF_buf4), );
  MUX2X1 MUX2X1_570 (.gnd(gnd), .A(_5394_), .Y(_5395_), .vdd(vdd), .B(_5383_), .S(_4033__bF_buf7), );
  OAI21X1 OAI21X1_2072 (.gnd(gnd), .A(_1663_), .Y(_5396_), .vdd(vdd), .B(raddr2_0_bF_buf83_), .C(raddr2_1_bF_buf0_), );
  AOI21X1 AOI21X1_356 (.gnd(gnd), .A(regs_16__29_), .Y(_5397_), .vdd(vdd), .B(raddr2_0_bF_buf82_), .C(_5396_), );
  NOR2X1 NOR2X1_242 (.gnd(gnd), .A(raddr2_0_bF_buf81_), .Y(_5398_), .vdd(vdd), .B(_1565_), );
  NAND2X1 NAND2X1_1071 (.gnd(gnd), .A(regs_18__29_), .Y(_5399_), .vdd(vdd), .B(raddr2_0_bF_buf80_), );
  NAND2X1 NAND2X1_1072 (.gnd(gnd), .A(_4038__bF_buf8), .Y(_5400_), .vdd(vdd), .B(_5399_), );
  OAI21X1 OAI21X1_2073 (.gnd(gnd), .A(_5400_), .Y(_5401_), .vdd(vdd), .B(_5398_), .C(raddr2_2_bF_buf8_), );
  OAI21X1 OAI21X1_2074 (.gnd(gnd), .A(_1466_), .Y(_5402_), .vdd(vdd), .B(raddr2_0_bF_buf79_), .C(raddr2_1_bF_buf14_bF_buf0_), );
  AOI21X1 AOI21X1_357 (.gnd(gnd), .A(regs_20__29_), .Y(_5403_), .vdd(vdd), .B(raddr2_0_bF_buf78_), .C(_5402_), );
  AND2X2 AND2X2_76 (.gnd(gnd), .A(regs_22__29_), .Y(_5404_), .vdd(vdd), .B(raddr2_0_bF_buf77_), );
  OAI21X1 OAI21X1_2075 (.gnd(gnd), .A(_1368_), .Y(_5405_), .vdd(vdd), .B(raddr2_0_bF_buf76_), .C(_4038__bF_buf7), );
  OAI21X1 OAI21X1_2076 (.gnd(gnd), .A(_5405_), .Y(_5406_), .vdd(vdd), .B(_5404_), .C(_4036__bF_buf3), );
  OAI22X1 OAI22X1_101 (.gnd(gnd), .A(_5397_), .Y(_5407_), .vdd(vdd), .B(_5401_), .C(_5406_), .D(_5403_), );
  NAND2X1 NAND2X1_1073 (.gnd(gnd), .A(regs_28__29_), .Y(_5408_), .vdd(vdd), .B(raddr2_0_bF_buf75_), );
  OAI21X1 OAI21X1_2077 (.gnd(gnd), .A(_3898_), .Y(_5409_), .vdd(vdd), .B(raddr2_0_bF_buf74_), .C(_5408_), );
  MUX2X1 MUX2X1_571 (.gnd(gnd), .A(_5409_), .Y(_5410_), .vdd(vdd), .B(regs_30__29_), .S(raddr2_1_bF_buf13_bF_buf0_), );
  NAND2X1 NAND2X1_1074 (.gnd(gnd), .A(regs_26__29_), .Y(_5411_), .vdd(vdd), .B(raddr2_0_bF_buf73_), );
  OAI21X1 OAI21X1_2078 (.gnd(gnd), .A(_1201_), .Y(_5412_), .vdd(vdd), .B(raddr2_0_bF_buf72_), .C(_5411_), );
  NAND2X1 NAND2X1_1075 (.gnd(gnd), .A(regs_24__29_), .Y(_5413_), .vdd(vdd), .B(raddr2_0_bF_buf71_), );
  OAI21X1 OAI21X1_2079 (.gnd(gnd), .A(_3895_), .Y(_5414_), .vdd(vdd), .B(raddr2_0_bF_buf70_), .C(_5413_), );
  MUX2X1 MUX2X1_572 (.gnd(gnd), .A(_5414_), .Y(_5415_), .vdd(vdd), .B(_5412_), .S(raddr2_1_bF_buf12_bF_buf0_), );
  MUX2X1 MUX2X1_573 (.gnd(gnd), .A(_5415_), .Y(_5416_), .vdd(vdd), .B(_5410_), .S(raddr2_2_bF_buf7_), );
  MUX2X1 MUX2X1_574 (.gnd(gnd), .A(_5416_), .Y(_5417_), .vdd(vdd), .B(_5407_), .S(_4033__bF_buf6), );
  MUX2X1 MUX2X1_575 (.gnd(gnd), .A(_5395_), .Y(_5512__29_), .vdd(vdd), .B(_5417_), .S(raddr2_4_bF_buf0_), );
  OAI21X1 OAI21X1_2080 (.gnd(gnd), .A(_3958_), .Y(_5418_), .vdd(vdd), .B(raddr2_0_bF_buf69_), .C(raddr2_1_bF_buf11_), );
  AOI21X1 AOI21X1_358 (.gnd(gnd), .A(regs_4__30_), .Y(_5419_), .vdd(vdd), .B(raddr2_0_bF_buf68_), .C(_5418_), );
  AND2X2 AND2X2_77 (.gnd(gnd), .A(regs_6__30_), .Y(_5420_), .vdd(vdd), .B(raddr2_0_bF_buf67_), );
  OAI21X1 OAI21X1_2081 (.gnd(gnd), .A(_2161_), .Y(_5421_), .vdd(vdd), .B(raddr2_0_bF_buf66_), .C(_4038__bF_buf6), );
  OAI21X1 OAI21X1_2082 (.gnd(gnd), .A(_5421_), .Y(_5422_), .vdd(vdd), .B(_5420_), .C(_4036__bF_buf2), );
  OAI21X1 OAI21X1_2083 (.gnd(gnd), .A(_3965_), .Y(_5423_), .vdd(vdd), .B(raddr2_0_bF_buf65_), .C(raddr2_1_bF_buf10_), );
  AOI21X1 AOI21X1_359 (.gnd(gnd), .A(regs_0__30_), .Y(_5424_), .vdd(vdd), .B(raddr2_0_bF_buf64_), .C(_5423_), );
  NOR2X1 NOR2X1_243 (.gnd(gnd), .A(raddr2_0_bF_buf63_), .Y(_5425_), .vdd(vdd), .B(_3962_), );
  NAND2X1 NAND2X1_1076 (.gnd(gnd), .A(regs_2__30_), .Y(_5426_), .vdd(vdd), .B(raddr2_0_bF_buf62_), );
  NAND2X1 NAND2X1_1077 (.gnd(gnd), .A(_4038__bF_buf5), .Y(_5427_), .vdd(vdd), .B(_5426_), );
  OAI21X1 OAI21X1_2084 (.gnd(gnd), .A(_5427_), .Y(_5428_), .vdd(vdd), .B(_5425_), .C(raddr2_2_bF_buf6_), );
  OAI22X1 OAI22X1_102 (.gnd(gnd), .A(_5424_), .Y(_5429_), .vdd(vdd), .B(_5428_), .C(_5422_), .D(_5419_), );
  NAND2X1 NAND2X1_1078 (.gnd(gnd), .A(regs_10__30_), .Y(_5430_), .vdd(vdd), .B(raddr2_0_bF_buf61_), );
  OAI21X1 OAI21X1_2085 (.gnd(gnd), .A(_1962_), .Y(_5431_), .vdd(vdd), .B(raddr2_0_bF_buf60_), .C(_5430_), );
  NAND2X1 NAND2X1_1079 (.gnd(gnd), .A(regs_8__30_), .Y(_5432_), .vdd(vdd), .B(raddr2_0_bF_buf59_), );
  OAI21X1 OAI21X1_2086 (.gnd(gnd), .A(_2060_), .Y(_5433_), .vdd(vdd), .B(raddr2_0_bF_buf58_), .C(_5432_), );
  MUX2X1 MUX2X1_576 (.gnd(gnd), .A(_5433_), .Y(_5434_), .vdd(vdd), .B(_5431_), .S(raddr2_1_bF_buf9_), );
  NAND2X1 NAND2X1_1080 (.gnd(gnd), .A(regs_14__30_), .Y(_5435_), .vdd(vdd), .B(raddr2_0_bF_buf57_), );
  OAI21X1 OAI21X1_2087 (.gnd(gnd), .A(_1765_), .Y(_5436_), .vdd(vdd), .B(raddr2_0_bF_buf56_), .C(_5435_), );
  NAND2X1 NAND2X1_1081 (.gnd(gnd), .A(regs_12__30_), .Y(_5437_), .vdd(vdd), .B(raddr2_0_bF_buf55_), );
  OAI21X1 OAI21X1_2088 (.gnd(gnd), .A(_1863_), .Y(_5438_), .vdd(vdd), .B(raddr2_0_bF_buf54_), .C(_5437_), );
  MUX2X1 MUX2X1_577 (.gnd(gnd), .A(_5438_), .Y(_5439_), .vdd(vdd), .B(_5436_), .S(raddr2_1_bF_buf8_), );
  MUX2X1 MUX2X1_578 (.gnd(gnd), .A(_5439_), .Y(_5440_), .vdd(vdd), .B(_5434_), .S(_4036__bF_buf1), );
  MUX2X1 MUX2X1_579 (.gnd(gnd), .A(_5440_), .Y(_5441_), .vdd(vdd), .B(_5429_), .S(_4033__bF_buf5), );
  OAI21X1 OAI21X1_2089 (.gnd(gnd), .A(_1665_), .Y(_5442_), .vdd(vdd), .B(raddr2_0_bF_buf53_), .C(raddr2_1_bF_buf7_), );
  AOI21X1 AOI21X1_360 (.gnd(gnd), .A(regs_16__30_), .Y(_5443_), .vdd(vdd), .B(raddr2_0_bF_buf52_), .C(_5442_), );
  NOR2X1 NOR2X1_244 (.gnd(gnd), .A(raddr2_0_bF_buf51_), .Y(_5444_), .vdd(vdd), .B(_1567_), );
  NAND2X1 NAND2X1_1082 (.gnd(gnd), .A(regs_18__30_), .Y(_5445_), .vdd(vdd), .B(raddr2_0_bF_buf50_), );
  NAND2X1 NAND2X1_1083 (.gnd(gnd), .A(_4038__bF_buf4), .Y(_5446_), .vdd(vdd), .B(_5445_), );
  OAI21X1 OAI21X1_2090 (.gnd(gnd), .A(_5446_), .Y(_5447_), .vdd(vdd), .B(_5444_), .C(raddr2_2_bF_buf5_), );
  OAI21X1 OAI21X1_2091 (.gnd(gnd), .A(_1468_), .Y(_5448_), .vdd(vdd), .B(raddr2_0_bF_buf49_), .C(raddr2_1_bF_buf6_), );
  AOI21X1 AOI21X1_361 (.gnd(gnd), .A(regs_20__30_), .Y(_5449_), .vdd(vdd), .B(raddr2_0_bF_buf48_), .C(_5448_), );
  AND2X2 AND2X2_78 (.gnd(gnd), .A(regs_22__30_), .Y(_5450_), .vdd(vdd), .B(raddr2_0_bF_buf47_), );
  OAI21X1 OAI21X1_2092 (.gnd(gnd), .A(_1370_), .Y(_5451_), .vdd(vdd), .B(raddr2_0_bF_buf46_), .C(_4038__bF_buf3), );
  OAI21X1 OAI21X1_2093 (.gnd(gnd), .A(_5451_), .Y(_5452_), .vdd(vdd), .B(_5450_), .C(_4036__bF_buf0), );
  OAI22X1 OAI22X1_103 (.gnd(gnd), .A(_5443_), .Y(_5453_), .vdd(vdd), .B(_5447_), .C(_5452_), .D(_5449_), );
  NAND2X1 NAND2X1_1084 (.gnd(gnd), .A(regs_28__30_), .Y(_5454_), .vdd(vdd), .B(raddr2_0_bF_buf45_), );
  OAI21X1 OAI21X1_2094 (.gnd(gnd), .A(_3944_), .Y(_5455_), .vdd(vdd), .B(raddr2_0_bF_buf44_), .C(_5454_), );
  MUX2X1 MUX2X1_580 (.gnd(gnd), .A(_5455_), .Y(_5456_), .vdd(vdd), .B(regs_30__30_), .S(raddr2_1_bF_buf5_), );
  NAND2X1 NAND2X1_1085 (.gnd(gnd), .A(regs_26__30_), .Y(_5457_), .vdd(vdd), .B(raddr2_0_bF_buf43_), );
  OAI21X1 OAI21X1_2095 (.gnd(gnd), .A(_1203_), .Y(_5458_), .vdd(vdd), .B(raddr2_0_bF_buf42_), .C(_5457_), );
  NAND2X1 NAND2X1_1086 (.gnd(gnd), .A(regs_24__30_), .Y(_5459_), .vdd(vdd), .B(raddr2_0_bF_buf41_), );
  OAI21X1 OAI21X1_2096 (.gnd(gnd), .A(_3950_), .Y(_5460_), .vdd(vdd), .B(raddr2_0_bF_buf40_), .C(_5459_), );
  MUX2X1 MUX2X1_581 (.gnd(gnd), .A(_5460_), .Y(_5461_), .vdd(vdd), .B(_5458_), .S(raddr2_1_bF_buf4_), );
  MUX2X1 MUX2X1_582 (.gnd(gnd), .A(_5461_), .Y(_5462_), .vdd(vdd), .B(_5456_), .S(raddr2_2_bF_buf4_), );
  MUX2X1 MUX2X1_583 (.gnd(gnd), .A(_5462_), .Y(_5463_), .vdd(vdd), .B(_5453_), .S(_4033__bF_buf4), );
  MUX2X1 MUX2X1_584 (.gnd(gnd), .A(_5441_), .Y(_5512__30_), .vdd(vdd), .B(_5463_), .S(raddr2_4_bF_buf4_), );
  NAND2X1 NAND2X1_1087 (.gnd(gnd), .A(regs_22__31_), .Y(_5464_), .vdd(vdd), .B(raddr2_0_bF_buf39_), );
  OAI21X1 OAI21X1_2097 (.gnd(gnd), .A(_1372_), .Y(_5465_), .vdd(vdd), .B(raddr2_0_bF_buf38_), .C(_5464_), );
  NAND2X1 NAND2X1_1088 (.gnd(gnd), .A(regs_20__31_), .Y(_5466_), .vdd(vdd), .B(raddr2_0_bF_buf37_), );
  OAI21X1 OAI21X1_2098 (.gnd(gnd), .A(_1470_), .Y(_5467_), .vdd(vdd), .B(raddr2_0_bF_buf36_), .C(_5466_), );
  MUX2X1 MUX2X1_585 (.gnd(gnd), .A(_5467_), .Y(_5468_), .vdd(vdd), .B(_5465_), .S(raddr2_1_bF_buf3_), );
  NAND2X1 NAND2X1_1089 (.gnd(gnd), .A(_4036__bF_buf8), .Y(_5469_), .vdd(vdd), .B(_5468_), );
  NAND2X1 NAND2X1_1090 (.gnd(gnd), .A(regs_18__31_), .Y(_5470_), .vdd(vdd), .B(raddr2_0_bF_buf35_), );
  OAI21X1 OAI21X1_2099 (.gnd(gnd), .A(_1569_), .Y(_5471_), .vdd(vdd), .B(raddr2_0_bF_buf34_), .C(_5470_), );
  NAND2X1 NAND2X1_1091 (.gnd(gnd), .A(regs_16__31_), .Y(_5472_), .vdd(vdd), .B(raddr2_0_bF_buf33_), );
  OAI21X1 OAI21X1_2100 (.gnd(gnd), .A(_1667_), .Y(_5473_), .vdd(vdd), .B(raddr2_0_bF_buf32_), .C(_5472_), );
  MUX2X1 MUX2X1_586 (.gnd(gnd), .A(_5473_), .Y(_5474_), .vdd(vdd), .B(_5471_), .S(raddr2_1_bF_buf2_), );
  AOI21X1 AOI21X1_362 (.gnd(gnd), .A(raddr2_2_bF_buf3_), .Y(_5475_), .vdd(vdd), .B(_5474_), .C(_4033__bF_buf3), );
  OAI21X1 OAI21X1_2101 (.gnd(gnd), .A(_1205_), .Y(_5476_), .vdd(vdd), .B(raddr2_0_bF_buf31_), .C(raddr2_2_bF_buf2_), );
  AOI21X1 AOI21X1_363 (.gnd(gnd), .A(regs_26__31_), .Y(_5477_), .vdd(vdd), .B(raddr2_0_bF_buf30_), .C(_5476_), );
  OAI21X1 OAI21X1_2102 (.gnd(gnd), .A(regs_30__31_), .Y(_5478_), .vdd(vdd), .B(raddr2_2_bF_buf1_), .C(_4038__bF_buf2), );
  OAI21X1 OAI21X1_2103 (.gnd(gnd), .A(_4027_), .Y(_5479_), .vdd(vdd), .B(raddr2_0_bF_buf29_), .C(raddr2_2_bF_buf0_), );
  AOI21X1 AOI21X1_364 (.gnd(gnd), .A(regs_24__31_), .Y(_5480_), .vdd(vdd), .B(raddr2_0_bF_buf28_), .C(_5479_), );
  NOR2X1 NOR2X1_245 (.gnd(gnd), .A(raddr2_0_bF_buf27_), .Y(_5481_), .vdd(vdd), .B(_4021_), );
  NAND2X1 NAND2X1_1092 (.gnd(gnd), .A(regs_28__31_), .Y(_5482_), .vdd(vdd), .B(raddr2_0_bF_buf26_), );
  NAND2X1 NAND2X1_1093 (.gnd(gnd), .A(_4036__bF_buf7), .Y(_5483_), .vdd(vdd), .B(_5482_), );
  OAI21X1 OAI21X1_2104 (.gnd(gnd), .A(_5483_), .Y(_5484_), .vdd(vdd), .B(_5481_), .C(raddr2_1_bF_buf1_), );
  OAI22X1 OAI22X1_104 (.gnd(gnd), .A(_5477_), .Y(_5485_), .vdd(vdd), .B(_5478_), .C(_5484_), .D(_5480_), );
  AOI22X1 AOI22X1_27 (.gnd(gnd), .A(_5485_), .Y(_5486_), .vdd(vdd), .B(_4033__bF_buf2), .C(_5469_), .D(_5475_), );
  OAI21X1 OAI21X1_2105 (.gnd(gnd), .A(_3982_), .Y(_5487_), .vdd(vdd), .B(raddr2_0_bF_buf25_), .C(raddr2_1_bF_buf0_), );
  AOI21X1 AOI21X1_365 (.gnd(gnd), .A(regs_4__31_), .Y(_5488_), .vdd(vdd), .B(raddr2_0_bF_buf24_), .C(_5487_), );
  AND2X2 AND2X2_79 (.gnd(gnd), .A(regs_6__31_), .Y(_5489_), .vdd(vdd), .B(raddr2_0_bF_buf23_), );
  OAI21X1 OAI21X1_2106 (.gnd(gnd), .A(_2163_), .Y(_5490_), .vdd(vdd), .B(raddr2_0_bF_buf22_), .C(_4038__bF_buf1), );
  OAI21X1 OAI21X1_2107 (.gnd(gnd), .A(_5490_), .Y(_5491_), .vdd(vdd), .B(_5489_), .C(_4036__bF_buf6), );
  OAI21X1 OAI21X1_2108 (.gnd(gnd), .A(_3988_), .Y(_5492_), .vdd(vdd), .B(raddr2_0_bF_buf21_), .C(raddr2_1_bF_buf14_bF_buf3_), );
  AOI21X1 AOI21X1_366 (.gnd(gnd), .A(regs_0__31_), .Y(_5493_), .vdd(vdd), .B(raddr2_0_bF_buf20_), .C(_5492_), );
  NOR2X1 NOR2X1_246 (.gnd(gnd), .A(raddr2_0_bF_buf19_), .Y(_5494_), .vdd(vdd), .B(_3991_), );
  NAND2X1 NAND2X1_1094 (.gnd(gnd), .A(regs_2__31_), .Y(_5495_), .vdd(vdd), .B(raddr2_0_bF_buf18_), );
  NAND2X1 NAND2X1_1095 (.gnd(gnd), .A(_4038__bF_buf0), .Y(_5496_), .vdd(vdd), .B(_5495_), );
  OAI21X1 OAI21X1_2109 (.gnd(gnd), .A(_5496_), .Y(_5497_), .vdd(vdd), .B(_5494_), .C(raddr2_2_bF_buf10_), );
  OAI22X1 OAI22X1_105 (.gnd(gnd), .A(_5493_), .Y(_5498_), .vdd(vdd), .B(_5497_), .C(_5491_), .D(_5488_), );
  NAND2X1 NAND2X1_1096 (.gnd(gnd), .A(regs_10__31_), .Y(_5499_), .vdd(vdd), .B(raddr2_0_bF_buf17_), );
  OAI21X1 OAI21X1_2110 (.gnd(gnd), .A(_1964_), .Y(_5500_), .vdd(vdd), .B(raddr2_0_bF_buf16_), .C(_5499_), );
  NAND2X1 NAND2X1_1097 (.gnd(gnd), .A(regs_8__31_), .Y(_5501_), .vdd(vdd), .B(raddr2_0_bF_buf15_), );
  OAI21X1 OAI21X1_2111 (.gnd(gnd), .A(_2062_), .Y(_5502_), .vdd(vdd), .B(raddr2_0_bF_buf14_), .C(_5501_), );
  MUX2X1 MUX2X1_587 (.gnd(gnd), .A(_5502_), .Y(_5503_), .vdd(vdd), .B(_5500_), .S(raddr2_1_bF_buf13_bF_buf3_), );
  NAND2X1 NAND2X1_1098 (.gnd(gnd), .A(regs_14__31_), .Y(_5504_), .vdd(vdd), .B(raddr2_0_bF_buf13_), );
  OAI21X1 OAI21X1_2112 (.gnd(gnd), .A(_1767_), .Y(_5505_), .vdd(vdd), .B(raddr2_0_bF_buf12_), .C(_5504_), );
  NAND2X1 NAND2X1_1099 (.gnd(gnd), .A(regs_12__31_), .Y(_5506_), .vdd(vdd), .B(raddr2_0_bF_buf11_), );
  OAI21X1 OAI21X1_2113 (.gnd(gnd), .A(_1865_), .Y(_5507_), .vdd(vdd), .B(raddr2_0_bF_buf10_), .C(_5506_), );
  MUX2X1 MUX2X1_588 (.gnd(gnd), .A(_5507_), .Y(_5508_), .vdd(vdd), .B(_5505_), .S(raddr2_1_bF_buf12_bF_buf3_), );
  MUX2X1 MUX2X1_589 (.gnd(gnd), .A(_5508_), .Y(_5509_), .vdd(vdd), .B(_5503_), .S(_4036__bF_buf5), );
  MUX2X1 MUX2X1_590 (.gnd(gnd), .A(_5509_), .Y(_5510_), .vdd(vdd), .B(_5498_), .S(_4033__bF_buf1), );
  MUX2X1 MUX2X1_591 (.gnd(gnd), .A(_5510_), .Y(_5512__31_), .vdd(vdd), .B(_5486_), .S(raddr2_4_bF_buf3_), );
  INVX8 INVX8_8 (.gnd(gnd), .A(wdata[0]), .Y(_992_), .vdd(vdd), );
  INVX1 INVX1_162 (.gnd(gnd), .A(waddr[4]), .Y(_993_), .vdd(vdd), );
  INVX1 INVX1_163 (.gnd(gnd), .A(waddr[3]), .Y(_994_), .vdd(vdd), );
  NAND2X1 NAND2X1_1100 (.gnd(gnd), .A(_993_), .Y(_995_), .vdd(vdd), .B(_994_), );
  NOR2X1 NOR2X1_247 (.gnd(gnd), .A(waddr[2]), .Y(_996_), .vdd(vdd), .B(_995_), );
  NAND2X1 NAND2X1_1101 (.gnd(gnd), .A(waddr[0]), .Y(_997_), .vdd(vdd), .B(wen), );
  NOR2X1 NOR2X1_248 (.gnd(gnd), .A(waddr[1]), .Y(_998_), .vdd(vdd), .B(_997_), );
  NAND2X1 NAND2X1_1102 (.gnd(gnd), .A(_998_), .Y(_999_), .vdd(vdd), .B(_996_), );
  INVX8 INVX8_9 (.gnd(gnd), .A(_996_), .Y(_1000_), .vdd(vdd), );
  INVX8 INVX8_10 (.gnd(gnd), .A(_998_), .Y(_1001_), .vdd(vdd), );
  OAI21X1 OAI21X1_2114 (.gnd(gnd), .A(_1000__bF_buf7), .Y(_1002_), .vdd(vdd), .B(_1001__bF_buf1), .C(regs_30__0_), );
  OAI21X1 OAI21X1_2115 (.gnd(gnd), .A(_992__bF_buf0), .Y(_736_), .vdd(vdd), .B(_999__bF_buf4), .C(_1002_), );
  INVX8 INVX8_11 (.gnd(gnd), .A(wdata[1]), .Y(_1003_), .vdd(vdd), );
  OAI21X1 OAI21X1_2116 (.gnd(gnd), .A(_1000__bF_buf6), .Y(_1004_), .vdd(vdd), .B(_1001__bF_buf0), .C(regs_30__1_), );
  OAI21X1 OAI21X1_2117 (.gnd(gnd), .A(_1003__bF_buf0), .Y(_747_), .vdd(vdd), .B(_999__bF_buf3), .C(_1004_), );
  INVX8 INVX8_12 (.gnd(gnd), .A(wdata[2]), .Y(_1005_), .vdd(vdd), );
  OAI21X1 OAI21X1_2118 (.gnd(gnd), .A(_1000__bF_buf5), .Y(_1006_), .vdd(vdd), .B(_1001__bF_buf9), .C(regs_30__2_), );
  OAI21X1 OAI21X1_2119 (.gnd(gnd), .A(_1005__bF_buf0), .Y(_758_), .vdd(vdd), .B(_999__bF_buf2), .C(_1006_), );
  INVX8 INVX8_13 (.gnd(gnd), .A(wdata[3]), .Y(_1007_), .vdd(vdd), );
  OAI21X1 OAI21X1_2120 (.gnd(gnd), .A(_1000__bF_buf4), .Y(_1008_), .vdd(vdd), .B(_1001__bF_buf8), .C(regs_30__3_), );
  OAI21X1 OAI21X1_2121 (.gnd(gnd), .A(_1007__bF_buf0), .Y(_761_), .vdd(vdd), .B(_999__bF_buf1), .C(_1008_), );
  INVX8 INVX8_14 (.gnd(gnd), .A(wdata[4]), .Y(_1009_), .vdd(vdd), );
  OAI21X1 OAI21X1_2122 (.gnd(gnd), .A(_1000__bF_buf3), .Y(_1010_), .vdd(vdd), .B(_1001__bF_buf7), .C(regs_30__4_), );
  OAI21X1 OAI21X1_2123 (.gnd(gnd), .A(_1009__bF_buf3), .Y(_762_), .vdd(vdd), .B(_999__bF_buf0), .C(_1010_), );
  INVX8 INVX8_15 (.gnd(gnd), .A(wdata[5]), .Y(_1011_), .vdd(vdd), );
  OAI21X1 OAI21X1_2124 (.gnd(gnd), .A(_1000__bF_buf2), .Y(_1012_), .vdd(vdd), .B(_1001__bF_buf6), .C(regs_30__5_), );
  OAI21X1 OAI21X1_2125 (.gnd(gnd), .A(_1011__bF_buf3), .Y(_763_), .vdd(vdd), .B(_999__bF_buf4), .C(_1012_), );
  INVX8 INVX8_16 (.gnd(gnd), .A(wdata[6]), .Y(_1013_), .vdd(vdd), );
  OAI21X1 OAI21X1_2126 (.gnd(gnd), .A(_1000__bF_buf1), .Y(_1014_), .vdd(vdd), .B(_1001__bF_buf5), .C(regs_30__6_), );
  OAI21X1 OAI21X1_2127 (.gnd(gnd), .A(_1013__bF_buf3), .Y(_764_), .vdd(vdd), .B(_999__bF_buf3), .C(_1014_), );
  INVX8 INVX8_17 (.gnd(gnd), .A(wdata[7]), .Y(_1015_), .vdd(vdd), );
  OAI21X1 OAI21X1_2128 (.gnd(gnd), .A(_1000__bF_buf0), .Y(_1016_), .vdd(vdd), .B(_1001__bF_buf4), .C(regs_30__7_), );
  OAI21X1 OAI21X1_2129 (.gnd(gnd), .A(_1015__bF_buf3), .Y(_765_), .vdd(vdd), .B(_999__bF_buf2), .C(_1016_), );
  INVX8 INVX8_18 (.gnd(gnd), .A(wdata[8]), .Y(_1017_), .vdd(vdd), );
  OAI21X1 OAI21X1_2130 (.gnd(gnd), .A(_1000__bF_buf7), .Y(_1018_), .vdd(vdd), .B(_1001__bF_buf3), .C(regs_30__8_), );
  OAI21X1 OAI21X1_2131 (.gnd(gnd), .A(_1017__bF_buf3), .Y(_766_), .vdd(vdd), .B(_999__bF_buf1), .C(_1018_), );
  INVX8 INVX8_19 (.gnd(gnd), .A(wdata[9]), .Y(_1019_), .vdd(vdd), );
  OAI21X1 OAI21X1_2132 (.gnd(gnd), .A(_1000__bF_buf6), .Y(_1020_), .vdd(vdd), .B(_1001__bF_buf2), .C(regs_30__9_), );
  OAI21X1 OAI21X1_2133 (.gnd(gnd), .A(_1019__bF_buf3), .Y(_767_), .vdd(vdd), .B(_999__bF_buf0), .C(_1020_), );
  INVX8 INVX8_20 (.gnd(gnd), .A(wdata[10]), .Y(_1021_), .vdd(vdd), );
  OAI21X1 OAI21X1_2134 (.gnd(gnd), .A(_1000__bF_buf5), .Y(_1022_), .vdd(vdd), .B(_1001__bF_buf1), .C(regs_30__10_), );
  OAI21X1 OAI21X1_2135 (.gnd(gnd), .A(_1021__bF_buf3), .Y(_737_), .vdd(vdd), .B(_999__bF_buf4), .C(_1022_), );
  INVX8 INVX8_21 (.gnd(gnd), .A(wdata[11]), .Y(_1023_), .vdd(vdd), );
  OAI21X1 OAI21X1_2136 (.gnd(gnd), .A(_1000__bF_buf4), .Y(_1024_), .vdd(vdd), .B(_1001__bF_buf0), .C(regs_30__11_), );
  OAI21X1 OAI21X1_2137 (.gnd(gnd), .A(_1023__bF_buf3), .Y(_738_), .vdd(vdd), .B(_999__bF_buf3), .C(_1024_), );
  INVX8 INVX8_22 (.gnd(gnd), .A(wdata[12]), .Y(_1025_), .vdd(vdd), );
  OAI21X1 OAI21X1_2138 (.gnd(gnd), .A(_1000__bF_buf3), .Y(_1026_), .vdd(vdd), .B(_1001__bF_buf9), .C(regs_30__12_), );
  OAI21X1 OAI21X1_2139 (.gnd(gnd), .A(_1025__bF_buf3), .Y(_739_), .vdd(vdd), .B(_999__bF_buf2), .C(_1026_), );
  INVX8 INVX8_23 (.gnd(gnd), .A(wdata[13]), .Y(_1027_), .vdd(vdd), );
  OAI21X1 OAI21X1_2140 (.gnd(gnd), .A(_1000__bF_buf2), .Y(_1028_), .vdd(vdd), .B(_1001__bF_buf8), .C(regs_30__13_), );
  OAI21X1 OAI21X1_2141 (.gnd(gnd), .A(_1027__bF_buf3), .Y(_740_), .vdd(vdd), .B(_999__bF_buf1), .C(_1028_), );
  INVX8 INVX8_24 (.gnd(gnd), .A(wdata[14]), .Y(_1029_), .vdd(vdd), );
  OAI21X1 OAI21X1_2142 (.gnd(gnd), .A(_1000__bF_buf1), .Y(_1030_), .vdd(vdd), .B(_1001__bF_buf7), .C(regs_30__14_), );
  OAI21X1 OAI21X1_2143 (.gnd(gnd), .A(_1029__bF_buf3), .Y(_741_), .vdd(vdd), .B(_999__bF_buf0), .C(_1030_), );
  INVX8 INVX8_25 (.gnd(gnd), .A(wdata[15]), .Y(_1031_), .vdd(vdd), );
  OAI21X1 OAI21X1_2144 (.gnd(gnd), .A(_1000__bF_buf0), .Y(_1032_), .vdd(vdd), .B(_1001__bF_buf6), .C(regs_30__15_), );
  OAI21X1 OAI21X1_2145 (.gnd(gnd), .A(_1031__bF_buf3), .Y(_742_), .vdd(vdd), .B(_999__bF_buf4), .C(_1032_), );
  INVX8 INVX8_26 (.gnd(gnd), .A(wdata[16]), .Y(_1033_), .vdd(vdd), );
  OAI21X1 OAI21X1_2146 (.gnd(gnd), .A(_1000__bF_buf7), .Y(_1034_), .vdd(vdd), .B(_1001__bF_buf5), .C(regs_30__16_), );
  OAI21X1 OAI21X1_2147 (.gnd(gnd), .A(_1033__bF_buf3), .Y(_743_), .vdd(vdd), .B(_999__bF_buf3), .C(_1034_), );
  INVX8 INVX8_27 (.gnd(gnd), .A(wdata[17]), .Y(_1035_), .vdd(vdd), );
  OAI21X1 OAI21X1_2148 (.gnd(gnd), .A(_1000__bF_buf6), .Y(_1036_), .vdd(vdd), .B(_1001__bF_buf4), .C(regs_30__17_), );
  OAI21X1 OAI21X1_2149 (.gnd(gnd), .A(_1035__bF_buf3), .Y(_744_), .vdd(vdd), .B(_999__bF_buf2), .C(_1036_), );
  INVX8 INVX8_28 (.gnd(gnd), .A(wdata[18]), .Y(_1037_), .vdd(vdd), );
  OAI21X1 OAI21X1_2150 (.gnd(gnd), .A(_1000__bF_buf5), .Y(_1038_), .vdd(vdd), .B(_1001__bF_buf3), .C(regs_30__18_), );
  OAI21X1 OAI21X1_2151 (.gnd(gnd), .A(_1037__bF_buf3), .Y(_745_), .vdd(vdd), .B(_999__bF_buf1), .C(_1038_), );
  INVX8 INVX8_29 (.gnd(gnd), .A(wdata[19]), .Y(_1039_), .vdd(vdd), );
  OAI21X1 OAI21X1_2152 (.gnd(gnd), .A(_1000__bF_buf4), .Y(_1040_), .vdd(vdd), .B(_1001__bF_buf2), .C(regs_30__19_), );
  OAI21X1 OAI21X1_2153 (.gnd(gnd), .A(_1039__bF_buf3), .Y(_746_), .vdd(vdd), .B(_999__bF_buf0), .C(_1040_), );
  INVX8 INVX8_30 (.gnd(gnd), .A(wdata[20]), .Y(_1041_), .vdd(vdd), );
  OAI21X1 OAI21X1_2154 (.gnd(gnd), .A(_1000__bF_buf3), .Y(_1042_), .vdd(vdd), .B(_1001__bF_buf1), .C(regs_30__20_), );
  OAI21X1 OAI21X1_2155 (.gnd(gnd), .A(_1041__bF_buf3), .Y(_748_), .vdd(vdd), .B(_999__bF_buf4), .C(_1042_), );
  INVX8 INVX8_31 (.gnd(gnd), .A(wdata[21]), .Y(_1043_), .vdd(vdd), );
  OAI21X1 OAI21X1_2156 (.gnd(gnd), .A(_1000__bF_buf2), .Y(_1044_), .vdd(vdd), .B(_1001__bF_buf0), .C(regs_30__21_), );
  OAI21X1 OAI21X1_2157 (.gnd(gnd), .A(_1043__bF_buf3), .Y(_749_), .vdd(vdd), .B(_999__bF_buf3), .C(_1044_), );
  INVX8 INVX8_32 (.gnd(gnd), .A(wdata[22]), .Y(_1045_), .vdd(vdd), );
  OAI21X1 OAI21X1_2158 (.gnd(gnd), .A(_1000__bF_buf1), .Y(_1046_), .vdd(vdd), .B(_1001__bF_buf9), .C(regs_30__22_), );
  OAI21X1 OAI21X1_2159 (.gnd(gnd), .A(_1045__bF_buf3), .Y(_750_), .vdd(vdd), .B(_999__bF_buf2), .C(_1046_), );
  INVX8 INVX8_33 (.gnd(gnd), .A(wdata[23]), .Y(_1047_), .vdd(vdd), );
  OAI21X1 OAI21X1_2160 (.gnd(gnd), .A(_1000__bF_buf0), .Y(_1048_), .vdd(vdd), .B(_1001__bF_buf8), .C(regs_30__23_), );
  OAI21X1 OAI21X1_2161 (.gnd(gnd), .A(_1047__bF_buf3), .Y(_751_), .vdd(vdd), .B(_999__bF_buf1), .C(_1048_), );
  INVX8 INVX8_34 (.gnd(gnd), .A(wdata[24]), .Y(_1049_), .vdd(vdd), );
  OAI21X1 OAI21X1_2162 (.gnd(gnd), .A(_1000__bF_buf7), .Y(_1050_), .vdd(vdd), .B(_1001__bF_buf7), .C(regs_30__24_), );
  OAI21X1 OAI21X1_2163 (.gnd(gnd), .A(_1049__bF_buf3), .Y(_752_), .vdd(vdd), .B(_999__bF_buf0), .C(_1050_), );
  INVX8 INVX8_35 (.gnd(gnd), .A(wdata[25]), .Y(_1051_), .vdd(vdd), );
  OAI21X1 OAI21X1_2164 (.gnd(gnd), .A(_1000__bF_buf6), .Y(_1052_), .vdd(vdd), .B(_1001__bF_buf6), .C(regs_30__25_), );
  OAI21X1 OAI21X1_2165 (.gnd(gnd), .A(_1051__bF_buf3), .Y(_753_), .vdd(vdd), .B(_999__bF_buf4), .C(_1052_), );
  INVX8 INVX8_36 (.gnd(gnd), .A(wdata[26]), .Y(_1053_), .vdd(vdd), );
  OAI21X1 OAI21X1_2166 (.gnd(gnd), .A(_1000__bF_buf5), .Y(_1054_), .vdd(vdd), .B(_1001__bF_buf5), .C(regs_30__26_), );
  OAI21X1 OAI21X1_2167 (.gnd(gnd), .A(_1053__bF_buf3), .Y(_754_), .vdd(vdd), .B(_999__bF_buf3), .C(_1054_), );
  INVX8 INVX8_37 (.gnd(gnd), .A(wdata[27]), .Y(_1055_), .vdd(vdd), );
  OAI21X1 OAI21X1_2168 (.gnd(gnd), .A(_1000__bF_buf4), .Y(_1056_), .vdd(vdd), .B(_1001__bF_buf4), .C(regs_30__27_), );
  OAI21X1 OAI21X1_2169 (.gnd(gnd), .A(_1055__bF_buf3), .Y(_755_), .vdd(vdd), .B(_999__bF_buf2), .C(_1056_), );
  INVX8 INVX8_38 (.gnd(gnd), .A(wdata[28]), .Y(_1057_), .vdd(vdd), );
  OAI21X1 OAI21X1_2170 (.gnd(gnd), .A(_1000__bF_buf3), .Y(_1058_), .vdd(vdd), .B(_1001__bF_buf3), .C(regs_30__28_), );
  OAI21X1 OAI21X1_2171 (.gnd(gnd), .A(_1057__bF_buf3), .Y(_756_), .vdd(vdd), .B(_999__bF_buf1), .C(_1058_), );
  INVX8 INVX8_39 (.gnd(gnd), .A(wdata[29]), .Y(_1059_), .vdd(vdd), );
  OAI21X1 OAI21X1_2172 (.gnd(gnd), .A(_1000__bF_buf2), .Y(_1060_), .vdd(vdd), .B(_1001__bF_buf2), .C(regs_30__29_), );
  OAI21X1 OAI21X1_2173 (.gnd(gnd), .A(_1059__bF_buf3), .Y(_757_), .vdd(vdd), .B(_999__bF_buf0), .C(_1060_), );
  INVX8 INVX8_40 (.gnd(gnd), .A(wdata[30]), .Y(_1061_), .vdd(vdd), );
  OAI21X1 OAI21X1_2174 (.gnd(gnd), .A(_1000__bF_buf1), .Y(_1062_), .vdd(vdd), .B(_1001__bF_buf1), .C(regs_30__30_), );
  OAI21X1 OAI21X1_2175 (.gnd(gnd), .A(_1061__bF_buf3), .Y(_759_), .vdd(vdd), .B(_999__bF_buf4), .C(_1062_), );
  INVX8 INVX8_41 (.gnd(gnd), .A(wdata[31]), .Y(_1063_), .vdd(vdd), );
  OAI21X1 OAI21X1_2176 (.gnd(gnd), .A(_1000__bF_buf0), .Y(_1064_), .vdd(vdd), .B(_1001__bF_buf0), .C(regs_30__31_), );
  OAI21X1 OAI21X1_2177 (.gnd(gnd), .A(_1063__bF_buf3), .Y(_760_), .vdd(vdd), .B(_999__bF_buf3), .C(_1064_), );
  INVX1 INVX1_164 (.gnd(gnd), .A(wen), .Y(_1065_), .vdd(vdd), );
  INVX1 INVX1_165 (.gnd(gnd), .A(waddr[0]), .Y(_1066_), .vdd(vdd), );
  NAND2X1 NAND2X1_1103 (.gnd(gnd), .A(waddr[1]), .Y(_1067_), .vdd(vdd), .B(_1066_), );
  NOR2X1 NOR2X1_249 (.gnd(gnd), .A(_1065_), .Y(_1068_), .vdd(vdd), .B(_1067_), );
  NAND2X1 NAND2X1_1104 (.gnd(gnd), .A(_1068_), .Y(_1069_), .vdd(vdd), .B(_996_), );
  INVX8 INVX8_42 (.gnd(gnd), .A(_1068_), .Y(_1070_), .vdd(vdd), );
  OAI21X1 OAI21X1_2178 (.gnd(gnd), .A(_1000__bF_buf7), .Y(_1071_), .vdd(vdd), .B(_1070__bF_buf8), .C(regs_29__0_), );
  OAI21X1 OAI21X1_2179 (.gnd(gnd), .A(_992__bF_buf3), .Y(_672_), .vdd(vdd), .B(_1069__bF_buf4), .C(_1071_), );
  OAI21X1 OAI21X1_2180 (.gnd(gnd), .A(_1000__bF_buf6), .Y(_1072_), .vdd(vdd), .B(_1070__bF_buf7), .C(regs_29__1_), );
  OAI21X1 OAI21X1_2181 (.gnd(gnd), .A(_1003__bF_buf3), .Y(_683_), .vdd(vdd), .B(_1069__bF_buf3), .C(_1072_), );
  OAI21X1 OAI21X1_2182 (.gnd(gnd), .A(_1000__bF_buf5), .Y(_1073_), .vdd(vdd), .B(_1070__bF_buf6), .C(regs_29__2_), );
  OAI21X1 OAI21X1_2183 (.gnd(gnd), .A(_1005__bF_buf3), .Y(_694_), .vdd(vdd), .B(_1069__bF_buf2), .C(_1073_), );
  OAI21X1 OAI21X1_2184 (.gnd(gnd), .A(_1000__bF_buf4), .Y(_1074_), .vdd(vdd), .B(_1070__bF_buf5), .C(regs_29__3_), );
  OAI21X1 OAI21X1_2185 (.gnd(gnd), .A(_1007__bF_buf3), .Y(_697_), .vdd(vdd), .B(_1069__bF_buf1), .C(_1074_), );
  OAI21X1 OAI21X1_2186 (.gnd(gnd), .A(_1000__bF_buf3), .Y(_1075_), .vdd(vdd), .B(_1070__bF_buf4), .C(regs_29__4_), );
  OAI21X1 OAI21X1_2187 (.gnd(gnd), .A(_1009__bF_buf2), .Y(_698_), .vdd(vdd), .B(_1069__bF_buf0), .C(_1075_), );
  OAI21X1 OAI21X1_2188 (.gnd(gnd), .A(_1000__bF_buf2), .Y(_1076_), .vdd(vdd), .B(_1070__bF_buf3), .C(regs_29__5_), );
  OAI21X1 OAI21X1_2189 (.gnd(gnd), .A(_1011__bF_buf2), .Y(_699_), .vdd(vdd), .B(_1069__bF_buf4), .C(_1076_), );
  OAI21X1 OAI21X1_2190 (.gnd(gnd), .A(_1000__bF_buf1), .Y(_1077_), .vdd(vdd), .B(_1070__bF_buf2), .C(regs_29__6_), );
  OAI21X1 OAI21X1_2191 (.gnd(gnd), .A(_1013__bF_buf2), .Y(_700_), .vdd(vdd), .B(_1069__bF_buf3), .C(_1077_), );
  OAI21X1 OAI21X1_2192 (.gnd(gnd), .A(_1000__bF_buf0), .Y(_1078_), .vdd(vdd), .B(_1070__bF_buf1), .C(regs_29__7_), );
  OAI21X1 OAI21X1_2193 (.gnd(gnd), .A(_1015__bF_buf2), .Y(_701_), .vdd(vdd), .B(_1069__bF_buf2), .C(_1078_), );
  OAI21X1 OAI21X1_2194 (.gnd(gnd), .A(_1000__bF_buf7), .Y(_1079_), .vdd(vdd), .B(_1070__bF_buf0), .C(regs_29__8_), );
  OAI21X1 OAI21X1_2195 (.gnd(gnd), .A(_1017__bF_buf2), .Y(_702_), .vdd(vdd), .B(_1069__bF_buf1), .C(_1079_), );
  OAI21X1 OAI21X1_2196 (.gnd(gnd), .A(_1000__bF_buf6), .Y(_1080_), .vdd(vdd), .B(_1070__bF_buf10), .C(regs_29__9_), );
  OAI21X1 OAI21X1_2197 (.gnd(gnd), .A(_1019__bF_buf2), .Y(_703_), .vdd(vdd), .B(_1069__bF_buf0), .C(_1080_), );
  OAI21X1 OAI21X1_2198 (.gnd(gnd), .A(_1000__bF_buf5), .Y(_1081_), .vdd(vdd), .B(_1070__bF_buf9), .C(regs_29__10_), );
  OAI21X1 OAI21X1_2199 (.gnd(gnd), .A(_1021__bF_buf2), .Y(_673_), .vdd(vdd), .B(_1069__bF_buf4), .C(_1081_), );
  OAI21X1 OAI21X1_2200 (.gnd(gnd), .A(_1000__bF_buf4), .Y(_1082_), .vdd(vdd), .B(_1070__bF_buf8), .C(regs_29__11_), );
  OAI21X1 OAI21X1_2201 (.gnd(gnd), .A(_1023__bF_buf2), .Y(_674_), .vdd(vdd), .B(_1069__bF_buf3), .C(_1082_), );
  OAI21X1 OAI21X1_2202 (.gnd(gnd), .A(_1000__bF_buf3), .Y(_1083_), .vdd(vdd), .B(_1070__bF_buf7), .C(regs_29__12_), );
  OAI21X1 OAI21X1_2203 (.gnd(gnd), .A(_1025__bF_buf2), .Y(_675_), .vdd(vdd), .B(_1069__bF_buf2), .C(_1083_), );
  OAI21X1 OAI21X1_2204 (.gnd(gnd), .A(_1000__bF_buf2), .Y(_1084_), .vdd(vdd), .B(_1070__bF_buf6), .C(regs_29__13_), );
  OAI21X1 OAI21X1_2205 (.gnd(gnd), .A(_1027__bF_buf2), .Y(_676_), .vdd(vdd), .B(_1069__bF_buf1), .C(_1084_), );
  OAI21X1 OAI21X1_2206 (.gnd(gnd), .A(_1000__bF_buf1), .Y(_1085_), .vdd(vdd), .B(_1070__bF_buf5), .C(regs_29__14_), );
  OAI21X1 OAI21X1_2207 (.gnd(gnd), .A(_1029__bF_buf2), .Y(_677_), .vdd(vdd), .B(_1069__bF_buf0), .C(_1085_), );
  OAI21X1 OAI21X1_2208 (.gnd(gnd), .A(_1000__bF_buf0), .Y(_1086_), .vdd(vdd), .B(_1070__bF_buf4), .C(regs_29__15_), );
  OAI21X1 OAI21X1_2209 (.gnd(gnd), .A(_1031__bF_buf2), .Y(_678_), .vdd(vdd), .B(_1069__bF_buf4), .C(_1086_), );
  OAI21X1 OAI21X1_2210 (.gnd(gnd), .A(_1000__bF_buf7), .Y(_1087_), .vdd(vdd), .B(_1070__bF_buf3), .C(regs_29__16_), );
  OAI21X1 OAI21X1_2211 (.gnd(gnd), .A(_1033__bF_buf2), .Y(_679_), .vdd(vdd), .B(_1069__bF_buf3), .C(_1087_), );
  OAI21X1 OAI21X1_2212 (.gnd(gnd), .A(_1000__bF_buf6), .Y(_1088_), .vdd(vdd), .B(_1070__bF_buf2), .C(regs_29__17_), );
  OAI21X1 OAI21X1_2213 (.gnd(gnd), .A(_1035__bF_buf2), .Y(_680_), .vdd(vdd), .B(_1069__bF_buf2), .C(_1088_), );
  OAI21X1 OAI21X1_2214 (.gnd(gnd), .A(_1000__bF_buf5), .Y(_1089_), .vdd(vdd), .B(_1070__bF_buf1), .C(regs_29__18_), );
  OAI21X1 OAI21X1_2215 (.gnd(gnd), .A(_1037__bF_buf2), .Y(_681_), .vdd(vdd), .B(_1069__bF_buf1), .C(_1089_), );
  OAI21X1 OAI21X1_2216 (.gnd(gnd), .A(_1000__bF_buf4), .Y(_1090_), .vdd(vdd), .B(_1070__bF_buf0), .C(regs_29__19_), );
  OAI21X1 OAI21X1_2217 (.gnd(gnd), .A(_1039__bF_buf2), .Y(_682_), .vdd(vdd), .B(_1069__bF_buf0), .C(_1090_), );
  OAI21X1 OAI21X1_2218 (.gnd(gnd), .A(_1000__bF_buf3), .Y(_1091_), .vdd(vdd), .B(_1070__bF_buf10), .C(regs_29__20_), );
  OAI21X1 OAI21X1_2219 (.gnd(gnd), .A(_1041__bF_buf2), .Y(_684_), .vdd(vdd), .B(_1069__bF_buf4), .C(_1091_), );
  OAI21X1 OAI21X1_2220 (.gnd(gnd), .A(_1000__bF_buf2), .Y(_1092_), .vdd(vdd), .B(_1070__bF_buf9), .C(regs_29__21_), );
  OAI21X1 OAI21X1_2221 (.gnd(gnd), .A(_1043__bF_buf2), .Y(_685_), .vdd(vdd), .B(_1069__bF_buf3), .C(_1092_), );
  OAI21X1 OAI21X1_2222 (.gnd(gnd), .A(_1000__bF_buf1), .Y(_1093_), .vdd(vdd), .B(_1070__bF_buf8), .C(regs_29__22_), );
  OAI21X1 OAI21X1_2223 (.gnd(gnd), .A(_1045__bF_buf2), .Y(_686_), .vdd(vdd), .B(_1069__bF_buf2), .C(_1093_), );
  OAI21X1 OAI21X1_2224 (.gnd(gnd), .A(_1000__bF_buf0), .Y(_1094_), .vdd(vdd), .B(_1070__bF_buf7), .C(regs_29__23_), );
  OAI21X1 OAI21X1_2225 (.gnd(gnd), .A(_1047__bF_buf2), .Y(_687_), .vdd(vdd), .B(_1069__bF_buf1), .C(_1094_), );
  OAI21X1 OAI21X1_2226 (.gnd(gnd), .A(_1000__bF_buf7), .Y(_1095_), .vdd(vdd), .B(_1070__bF_buf6), .C(regs_29__24_), );
  OAI21X1 OAI21X1_2227 (.gnd(gnd), .A(_1049__bF_buf2), .Y(_688_), .vdd(vdd), .B(_1069__bF_buf0), .C(_1095_), );
  OAI21X1 OAI21X1_2228 (.gnd(gnd), .A(_1000__bF_buf6), .Y(_1096_), .vdd(vdd), .B(_1070__bF_buf5), .C(regs_29__25_), );
  OAI21X1 OAI21X1_2229 (.gnd(gnd), .A(_1051__bF_buf2), .Y(_689_), .vdd(vdd), .B(_1069__bF_buf4), .C(_1096_), );
  OAI21X1 OAI21X1_2230 (.gnd(gnd), .A(_1000__bF_buf5), .Y(_1097_), .vdd(vdd), .B(_1070__bF_buf4), .C(regs_29__26_), );
  OAI21X1 OAI21X1_2231 (.gnd(gnd), .A(_1053__bF_buf2), .Y(_690_), .vdd(vdd), .B(_1069__bF_buf3), .C(_1097_), );
  OAI21X1 OAI21X1_2232 (.gnd(gnd), .A(_1000__bF_buf4), .Y(_1098_), .vdd(vdd), .B(_1070__bF_buf3), .C(regs_29__27_), );
  OAI21X1 OAI21X1_2233 (.gnd(gnd), .A(_1055__bF_buf2), .Y(_691_), .vdd(vdd), .B(_1069__bF_buf2), .C(_1098_), );
  OAI21X1 OAI21X1_2234 (.gnd(gnd), .A(_1000__bF_buf3), .Y(_1099_), .vdd(vdd), .B(_1070__bF_buf2), .C(regs_29__28_), );
  OAI21X1 OAI21X1_2235 (.gnd(gnd), .A(_1057__bF_buf2), .Y(_692_), .vdd(vdd), .B(_1069__bF_buf1), .C(_1099_), );
  OAI21X1 OAI21X1_2236 (.gnd(gnd), .A(_1000__bF_buf2), .Y(_1100_), .vdd(vdd), .B(_1070__bF_buf1), .C(regs_29__29_), );
  OAI21X1 OAI21X1_2237 (.gnd(gnd), .A(_1059__bF_buf2), .Y(_693_), .vdd(vdd), .B(_1069__bF_buf0), .C(_1100_), );
  OAI21X1 OAI21X1_2238 (.gnd(gnd), .A(_1000__bF_buf1), .Y(_1101_), .vdd(vdd), .B(_1070__bF_buf0), .C(regs_29__30_), );
  OAI21X1 OAI21X1_2239 (.gnd(gnd), .A(_1061__bF_buf2), .Y(_695_), .vdd(vdd), .B(_1069__bF_buf4), .C(_1101_), );
  OAI21X1 OAI21X1_2240 (.gnd(gnd), .A(_1000__bF_buf0), .Y(_1102_), .vdd(vdd), .B(_1070__bF_buf10), .C(regs_29__31_), );
  OAI21X1 OAI21X1_2241 (.gnd(gnd), .A(_1063__bF_buf2), .Y(_696_), .vdd(vdd), .B(_1069__bF_buf3), .C(_1102_), );
  INVX1 INVX1_166 (.gnd(gnd), .A(waddr[1]), .Y(_1103_), .vdd(vdd), );
  OR2X2 OR2X2_11 (.gnd(gnd), .A(_997_), .Y(_1104_), .vdd(vdd), .B(_1103_), );
  NOR2X1 NOR2X1_250 (.gnd(gnd), .A(_1104__bF_buf0), .Y(_1105_), .vdd(vdd), .B(_1000__bF_buf7), );
  NOR2X1 NOR2X1_251 (.gnd(gnd), .A(regs_28__0_), .Y(_1106_), .vdd(vdd), .B(_1105__bF_buf7), );
  AOI21X1 AOI21X1_367 (.gnd(gnd), .A(_992__bF_buf2), .Y(_640_), .vdd(vdd), .B(_1105__bF_buf6), .C(_1106_), );
  NOR2X1 NOR2X1_252 (.gnd(gnd), .A(regs_28__1_), .Y(_1107_), .vdd(vdd), .B(_1105__bF_buf5), );
  AOI21X1 AOI21X1_368 (.gnd(gnd), .A(_1003__bF_buf2), .Y(_651_), .vdd(vdd), .B(_1105__bF_buf4), .C(_1107_), );
  NOR2X1 NOR2X1_253 (.gnd(gnd), .A(regs_28__2_), .Y(_1108_), .vdd(vdd), .B(_1105__bF_buf3), );
  AOI21X1 AOI21X1_369 (.gnd(gnd), .A(_1005__bF_buf2), .Y(_662_), .vdd(vdd), .B(_1105__bF_buf2), .C(_1108_), );
  NOR2X1 NOR2X1_254 (.gnd(gnd), .A(regs_28__3_), .Y(_1109_), .vdd(vdd), .B(_1105__bF_buf1), );
  AOI21X1 AOI21X1_370 (.gnd(gnd), .A(_1007__bF_buf2), .Y(_665_), .vdd(vdd), .B(_1105__bF_buf0), .C(_1109_), );
  NOR2X1 NOR2X1_255 (.gnd(gnd), .A(regs_28__4_), .Y(_1110_), .vdd(vdd), .B(_1105__bF_buf7), );
  AOI21X1 AOI21X1_371 (.gnd(gnd), .A(_1009__bF_buf1), .Y(_666_), .vdd(vdd), .B(_1105__bF_buf6), .C(_1110_), );
  NOR2X1 NOR2X1_256 (.gnd(gnd), .A(regs_28__5_), .Y(_1111_), .vdd(vdd), .B(_1105__bF_buf5), );
  AOI21X1 AOI21X1_372 (.gnd(gnd), .A(_1011__bF_buf1), .Y(_667_), .vdd(vdd), .B(_1105__bF_buf4), .C(_1111_), );
  NOR2X1 NOR2X1_257 (.gnd(gnd), .A(regs_28__6_), .Y(_1112_), .vdd(vdd), .B(_1105__bF_buf3), );
  AOI21X1 AOI21X1_373 (.gnd(gnd), .A(_1013__bF_buf1), .Y(_668_), .vdd(vdd), .B(_1105__bF_buf2), .C(_1112_), );
  NOR2X1 NOR2X1_258 (.gnd(gnd), .A(regs_28__7_), .Y(_1113_), .vdd(vdd), .B(_1105__bF_buf1), );
  AOI21X1 AOI21X1_374 (.gnd(gnd), .A(_1015__bF_buf1), .Y(_669_), .vdd(vdd), .B(_1105__bF_buf0), .C(_1113_), );
  NOR2X1 NOR2X1_259 (.gnd(gnd), .A(regs_28__8_), .Y(_1114_), .vdd(vdd), .B(_1105__bF_buf7), );
  AOI21X1 AOI21X1_375 (.gnd(gnd), .A(_1017__bF_buf1), .Y(_670_), .vdd(vdd), .B(_1105__bF_buf6), .C(_1114_), );
  NOR2X1 NOR2X1_260 (.gnd(gnd), .A(regs_28__9_), .Y(_1115_), .vdd(vdd), .B(_1105__bF_buf5), );
  AOI21X1 AOI21X1_376 (.gnd(gnd), .A(_1019__bF_buf1), .Y(_671_), .vdd(vdd), .B(_1105__bF_buf4), .C(_1115_), );
  NOR2X1 NOR2X1_261 (.gnd(gnd), .A(regs_28__10_), .Y(_1116_), .vdd(vdd), .B(_1105__bF_buf3), );
  AOI21X1 AOI21X1_377 (.gnd(gnd), .A(_1021__bF_buf1), .Y(_641_), .vdd(vdd), .B(_1105__bF_buf2), .C(_1116_), );
  NOR2X1 NOR2X1_262 (.gnd(gnd), .A(regs_28__11_), .Y(_1117_), .vdd(vdd), .B(_1105__bF_buf1), );
  AOI21X1 AOI21X1_378 (.gnd(gnd), .A(_1023__bF_buf1), .Y(_642_), .vdd(vdd), .B(_1105__bF_buf0), .C(_1117_), );
  NOR2X1 NOR2X1_263 (.gnd(gnd), .A(regs_28__12_), .Y(_1118_), .vdd(vdd), .B(_1105__bF_buf7), );
  AOI21X1 AOI21X1_379 (.gnd(gnd), .A(_1025__bF_buf1), .Y(_643_), .vdd(vdd), .B(_1105__bF_buf6), .C(_1118_), );
  NOR2X1 NOR2X1_264 (.gnd(gnd), .A(regs_28__13_), .Y(_1119_), .vdd(vdd), .B(_1105__bF_buf5), );
  AOI21X1 AOI21X1_380 (.gnd(gnd), .A(_1027__bF_buf1), .Y(_644_), .vdd(vdd), .B(_1105__bF_buf4), .C(_1119_), );
  NOR2X1 NOR2X1_265 (.gnd(gnd), .A(regs_28__14_), .Y(_1120_), .vdd(vdd), .B(_1105__bF_buf3), );
  AOI21X1 AOI21X1_381 (.gnd(gnd), .A(_1029__bF_buf1), .Y(_645_), .vdd(vdd), .B(_1105__bF_buf2), .C(_1120_), );
  NOR2X1 NOR2X1_266 (.gnd(gnd), .A(regs_28__15_), .Y(_1121_), .vdd(vdd), .B(_1105__bF_buf1), );
  AOI21X1 AOI21X1_382 (.gnd(gnd), .A(_1031__bF_buf1), .Y(_646_), .vdd(vdd), .B(_1105__bF_buf0), .C(_1121_), );
  NOR2X1 NOR2X1_267 (.gnd(gnd), .A(regs_28__16_), .Y(_1122_), .vdd(vdd), .B(_1105__bF_buf7), );
  AOI21X1 AOI21X1_383 (.gnd(gnd), .A(_1033__bF_buf1), .Y(_647_), .vdd(vdd), .B(_1105__bF_buf6), .C(_1122_), );
  NOR2X1 NOR2X1_268 (.gnd(gnd), .A(regs_28__17_), .Y(_1123_), .vdd(vdd), .B(_1105__bF_buf5), );
  AOI21X1 AOI21X1_384 (.gnd(gnd), .A(_1035__bF_buf1), .Y(_648_), .vdd(vdd), .B(_1105__bF_buf4), .C(_1123_), );
  NOR2X1 NOR2X1_269 (.gnd(gnd), .A(regs_28__18_), .Y(_1124_), .vdd(vdd), .B(_1105__bF_buf3), );
  AOI21X1 AOI21X1_385 (.gnd(gnd), .A(_1037__bF_buf1), .Y(_649_), .vdd(vdd), .B(_1105__bF_buf2), .C(_1124_), );
  NOR2X1 NOR2X1_270 (.gnd(gnd), .A(regs_28__19_), .Y(_1125_), .vdd(vdd), .B(_1105__bF_buf1), );
  AOI21X1 AOI21X1_386 (.gnd(gnd), .A(_1039__bF_buf1), .Y(_650_), .vdd(vdd), .B(_1105__bF_buf0), .C(_1125_), );
  NOR2X1 NOR2X1_271 (.gnd(gnd), .A(regs_28__20_), .Y(_1126_), .vdd(vdd), .B(_1105__bF_buf7), );
  AOI21X1 AOI21X1_387 (.gnd(gnd), .A(_1041__bF_buf1), .Y(_652_), .vdd(vdd), .B(_1105__bF_buf6), .C(_1126_), );
  NOR2X1 NOR2X1_272 (.gnd(gnd), .A(regs_28__21_), .Y(_1127_), .vdd(vdd), .B(_1105__bF_buf5), );
  AOI21X1 AOI21X1_388 (.gnd(gnd), .A(_1043__bF_buf1), .Y(_653_), .vdd(vdd), .B(_1105__bF_buf4), .C(_1127_), );
  NOR2X1 NOR2X1_273 (.gnd(gnd), .A(regs_28__22_), .Y(_1128_), .vdd(vdd), .B(_1105__bF_buf3), );
  AOI21X1 AOI21X1_389 (.gnd(gnd), .A(_1045__bF_buf1), .Y(_654_), .vdd(vdd), .B(_1105__bF_buf2), .C(_1128_), );
  NOR2X1 NOR2X1_274 (.gnd(gnd), .A(regs_28__23_), .Y(_1129_), .vdd(vdd), .B(_1105__bF_buf1), );
  AOI21X1 AOI21X1_390 (.gnd(gnd), .A(_1047__bF_buf1), .Y(_655_), .vdd(vdd), .B(_1105__bF_buf0), .C(_1129_), );
  NOR2X1 NOR2X1_275 (.gnd(gnd), .A(regs_28__24_), .Y(_1130_), .vdd(vdd), .B(_1105__bF_buf7), );
  AOI21X1 AOI21X1_391 (.gnd(gnd), .A(_1049__bF_buf1), .Y(_656_), .vdd(vdd), .B(_1105__bF_buf6), .C(_1130_), );
  NOR2X1 NOR2X1_276 (.gnd(gnd), .A(regs_28__25_), .Y(_1131_), .vdd(vdd), .B(_1105__bF_buf5), );
  AOI21X1 AOI21X1_392 (.gnd(gnd), .A(_1051__bF_buf1), .Y(_657_), .vdd(vdd), .B(_1105__bF_buf4), .C(_1131_), );
  NOR2X1 NOR2X1_277 (.gnd(gnd), .A(regs_28__26_), .Y(_1132_), .vdd(vdd), .B(_1105__bF_buf3), );
  AOI21X1 AOI21X1_393 (.gnd(gnd), .A(_1053__bF_buf1), .Y(_658_), .vdd(vdd), .B(_1105__bF_buf2), .C(_1132_), );
  NOR2X1 NOR2X1_278 (.gnd(gnd), .A(regs_28__27_), .Y(_1133_), .vdd(vdd), .B(_1105__bF_buf1), );
  AOI21X1 AOI21X1_394 (.gnd(gnd), .A(_1055__bF_buf1), .Y(_659_), .vdd(vdd), .B(_1105__bF_buf0), .C(_1133_), );
  NOR2X1 NOR2X1_279 (.gnd(gnd), .A(regs_28__28_), .Y(_1134_), .vdd(vdd), .B(_1105__bF_buf7), );
  AOI21X1 AOI21X1_395 (.gnd(gnd), .A(_1057__bF_buf1), .Y(_660_), .vdd(vdd), .B(_1105__bF_buf6), .C(_1134_), );
  NOR2X1 NOR2X1_280 (.gnd(gnd), .A(regs_28__29_), .Y(_1135_), .vdd(vdd), .B(_1105__bF_buf5), );
  AOI21X1 AOI21X1_396 (.gnd(gnd), .A(_1059__bF_buf1), .Y(_661_), .vdd(vdd), .B(_1105__bF_buf4), .C(_1135_), );
  NOR2X1 NOR2X1_281 (.gnd(gnd), .A(regs_28__30_), .Y(_1136_), .vdd(vdd), .B(_1105__bF_buf3), );
  AOI21X1 AOI21X1_397 (.gnd(gnd), .A(_1061__bF_buf1), .Y(_663_), .vdd(vdd), .B(_1105__bF_buf2), .C(_1136_), );
  NOR2X1 NOR2X1_282 (.gnd(gnd), .A(regs_28__31_), .Y(_1137_), .vdd(vdd), .B(_1105__bF_buf1), );
  AOI21X1 AOI21X1_398 (.gnd(gnd), .A(_1063__bF_buf1), .Y(_664_), .vdd(vdd), .B(_1105__bF_buf0), .C(_1137_), );
  INVX2 INVX2_289 (.gnd(gnd), .A(regs_27__0_), .Y(_1138_), .vdd(vdd), );
  INVX2 INVX2_290 (.gnd(gnd), .A(waddr[2]), .Y(_1139_), .vdd(vdd), );
  NOR2X1 NOR2X1_283 (.gnd(gnd), .A(_1139_), .Y(_1140_), .vdd(vdd), .B(_995_), );
  INVX8 INVX8_43 (.gnd(gnd), .A(_1140_), .Y(_1141_), .vdd(vdd), );
  NAND3X1 NAND3X1_1 (.gnd(gnd), .A(wen), .Y(_1142_), .vdd(vdd), .B(_1103_), .C(_1066_), );
  NOR2X1 NOR2X1_284 (.gnd(gnd), .A(_1142__bF_buf3), .Y(_1143_), .vdd(vdd), .B(_1141__bF_buf3), );
  NAND2X1 NAND2X1_1105 (.gnd(gnd), .A(wdata[0]), .Y(_1144_), .vdd(vdd), .B(_1143__bF_buf7), );
  OAI21X1 OAI21X1_2242 (.gnd(gnd), .A(_1138_), .Y(_608_), .vdd(vdd), .B(_1143__bF_buf6), .C(_1144_), );
  INVX2 INVX2_291 (.gnd(gnd), .A(regs_27__1_), .Y(_1145_), .vdd(vdd), );
  NAND2X1 NAND2X1_1106 (.gnd(gnd), .A(wdata[1]), .Y(_1146_), .vdd(vdd), .B(_1143__bF_buf5), );
  OAI21X1 OAI21X1_2243 (.gnd(gnd), .A(_1145_), .Y(_619_), .vdd(vdd), .B(_1143__bF_buf4), .C(_1146_), );
  INVX2 INVX2_292 (.gnd(gnd), .A(regs_27__2_), .Y(_1147_), .vdd(vdd), );
  NAND2X1 NAND2X1_1107 (.gnd(gnd), .A(wdata[2]), .Y(_1148_), .vdd(vdd), .B(_1143__bF_buf3), );
  OAI21X1 OAI21X1_2244 (.gnd(gnd), .A(_1147_), .Y(_630_), .vdd(vdd), .B(_1143__bF_buf2), .C(_1148_), );
  INVX2 INVX2_293 (.gnd(gnd), .A(regs_27__3_), .Y(_1149_), .vdd(vdd), );
  NAND2X1 NAND2X1_1108 (.gnd(gnd), .A(wdata[3]), .Y(_1150_), .vdd(vdd), .B(_1143__bF_buf1), );
  OAI21X1 OAI21X1_2245 (.gnd(gnd), .A(_1149_), .Y(_633_), .vdd(vdd), .B(_1143__bF_buf0), .C(_1150_), );
  INVX2 INVX2_294 (.gnd(gnd), .A(regs_27__4_), .Y(_1151_), .vdd(vdd), );
  NAND2X1 NAND2X1_1109 (.gnd(gnd), .A(wdata[4]), .Y(_1152_), .vdd(vdd), .B(_1143__bF_buf7), );
  OAI21X1 OAI21X1_2246 (.gnd(gnd), .A(_1151_), .Y(_634_), .vdd(vdd), .B(_1143__bF_buf6), .C(_1152_), );
  INVX2 INVX2_295 (.gnd(gnd), .A(regs_27__5_), .Y(_1153_), .vdd(vdd), );
  NAND2X1 NAND2X1_1110 (.gnd(gnd), .A(wdata[5]), .Y(_1154_), .vdd(vdd), .B(_1143__bF_buf5), );
  OAI21X1 OAI21X1_2247 (.gnd(gnd), .A(_1153_), .Y(_635_), .vdd(vdd), .B(_1143__bF_buf4), .C(_1154_), );
  INVX2 INVX2_296 (.gnd(gnd), .A(regs_27__6_), .Y(_1155_), .vdd(vdd), );
  NAND2X1 NAND2X1_1111 (.gnd(gnd), .A(wdata[6]), .Y(_1156_), .vdd(vdd), .B(_1143__bF_buf3), );
  OAI21X1 OAI21X1_2248 (.gnd(gnd), .A(_1155_), .Y(_636_), .vdd(vdd), .B(_1143__bF_buf2), .C(_1156_), );
  INVX2 INVX2_297 (.gnd(gnd), .A(regs_27__7_), .Y(_1157_), .vdd(vdd), );
  NAND2X1 NAND2X1_1112 (.gnd(gnd), .A(wdata[7]), .Y(_1158_), .vdd(vdd), .B(_1143__bF_buf1), );
  OAI21X1 OAI21X1_2249 (.gnd(gnd), .A(_1157_), .Y(_637_), .vdd(vdd), .B(_1143__bF_buf0), .C(_1158_), );
  INVX2 INVX2_298 (.gnd(gnd), .A(regs_27__8_), .Y(_1159_), .vdd(vdd), );
  NAND2X1 NAND2X1_1113 (.gnd(gnd), .A(wdata[8]), .Y(_1160_), .vdd(vdd), .B(_1143__bF_buf7), );
  OAI21X1 OAI21X1_2250 (.gnd(gnd), .A(_1159_), .Y(_638_), .vdd(vdd), .B(_1143__bF_buf6), .C(_1160_), );
  INVX2 INVX2_299 (.gnd(gnd), .A(regs_27__9_), .Y(_1161_), .vdd(vdd), );
  NAND2X1 NAND2X1_1114 (.gnd(gnd), .A(wdata[9]), .Y(_1162_), .vdd(vdd), .B(_1143__bF_buf5), );
  OAI21X1 OAI21X1_2251 (.gnd(gnd), .A(_1161_), .Y(_639_), .vdd(vdd), .B(_1143__bF_buf4), .C(_1162_), );
  INVX2 INVX2_300 (.gnd(gnd), .A(regs_27__10_), .Y(_1163_), .vdd(vdd), );
  NAND2X1 NAND2X1_1115 (.gnd(gnd), .A(wdata[10]), .Y(_1164_), .vdd(vdd), .B(_1143__bF_buf3), );
  OAI21X1 OAI21X1_2252 (.gnd(gnd), .A(_1163_), .Y(_609_), .vdd(vdd), .B(_1143__bF_buf2), .C(_1164_), );
  INVX2 INVX2_301 (.gnd(gnd), .A(regs_27__11_), .Y(_1165_), .vdd(vdd), );
  NAND2X1 NAND2X1_1116 (.gnd(gnd), .A(wdata[11]), .Y(_1166_), .vdd(vdd), .B(_1143__bF_buf1), );
  OAI21X1 OAI21X1_2253 (.gnd(gnd), .A(_1165_), .Y(_610_), .vdd(vdd), .B(_1143__bF_buf0), .C(_1166_), );
  INVX2 INVX2_302 (.gnd(gnd), .A(regs_27__12_), .Y(_1167_), .vdd(vdd), );
  NAND2X1 NAND2X1_1117 (.gnd(gnd), .A(wdata[12]), .Y(_1168_), .vdd(vdd), .B(_1143__bF_buf7), );
  OAI21X1 OAI21X1_2254 (.gnd(gnd), .A(_1167_), .Y(_611_), .vdd(vdd), .B(_1143__bF_buf6), .C(_1168_), );
  INVX2 INVX2_303 (.gnd(gnd), .A(regs_27__13_), .Y(_1169_), .vdd(vdd), );
  NAND2X1 NAND2X1_1118 (.gnd(gnd), .A(wdata[13]), .Y(_1170_), .vdd(vdd), .B(_1143__bF_buf5), );
  OAI21X1 OAI21X1_2255 (.gnd(gnd), .A(_1169_), .Y(_612_), .vdd(vdd), .B(_1143__bF_buf4), .C(_1170_), );
  INVX2 INVX2_304 (.gnd(gnd), .A(regs_27__14_), .Y(_1171_), .vdd(vdd), );
  NAND2X1 NAND2X1_1119 (.gnd(gnd), .A(wdata[14]), .Y(_1172_), .vdd(vdd), .B(_1143__bF_buf3), );
  OAI21X1 OAI21X1_2256 (.gnd(gnd), .A(_1171_), .Y(_613_), .vdd(vdd), .B(_1143__bF_buf2), .C(_1172_), );
  INVX2 INVX2_305 (.gnd(gnd), .A(regs_27__15_), .Y(_1173_), .vdd(vdd), );
  NAND2X1 NAND2X1_1120 (.gnd(gnd), .A(wdata[15]), .Y(_1174_), .vdd(vdd), .B(_1143__bF_buf1), );
  OAI21X1 OAI21X1_2257 (.gnd(gnd), .A(_1173_), .Y(_614_), .vdd(vdd), .B(_1143__bF_buf0), .C(_1174_), );
  INVX2 INVX2_306 (.gnd(gnd), .A(regs_27__16_), .Y(_1175_), .vdd(vdd), );
  NAND2X1 NAND2X1_1121 (.gnd(gnd), .A(wdata[16]), .Y(_1176_), .vdd(vdd), .B(_1143__bF_buf7), );
  OAI21X1 OAI21X1_2258 (.gnd(gnd), .A(_1175_), .Y(_615_), .vdd(vdd), .B(_1143__bF_buf6), .C(_1176_), );
  INVX2 INVX2_307 (.gnd(gnd), .A(regs_27__17_), .Y(_1177_), .vdd(vdd), );
  NAND2X1 NAND2X1_1122 (.gnd(gnd), .A(wdata[17]), .Y(_1178_), .vdd(vdd), .B(_1143__bF_buf5), );
  OAI21X1 OAI21X1_2259 (.gnd(gnd), .A(_1177_), .Y(_616_), .vdd(vdd), .B(_1143__bF_buf4), .C(_1178_), );
  INVX2 INVX2_308 (.gnd(gnd), .A(regs_27__18_), .Y(_1179_), .vdd(vdd), );
  NAND2X1 NAND2X1_1123 (.gnd(gnd), .A(wdata[18]), .Y(_1180_), .vdd(vdd), .B(_1143__bF_buf3), );
  OAI21X1 OAI21X1_2260 (.gnd(gnd), .A(_1179_), .Y(_617_), .vdd(vdd), .B(_1143__bF_buf2), .C(_1180_), );
  INVX2 INVX2_309 (.gnd(gnd), .A(regs_27__19_), .Y(_1181_), .vdd(vdd), );
  NAND2X1 NAND2X1_1124 (.gnd(gnd), .A(wdata[19]), .Y(_1182_), .vdd(vdd), .B(_1143__bF_buf1), );
  OAI21X1 OAI21X1_2261 (.gnd(gnd), .A(_1181_), .Y(_618_), .vdd(vdd), .B(_1143__bF_buf0), .C(_1182_), );
  INVX2 INVX2_310 (.gnd(gnd), .A(regs_27__20_), .Y(_1183_), .vdd(vdd), );
  NAND2X1 NAND2X1_1125 (.gnd(gnd), .A(wdata[20]), .Y(_1184_), .vdd(vdd), .B(_1143__bF_buf7), );
  OAI21X1 OAI21X1_2262 (.gnd(gnd), .A(_1183_), .Y(_620_), .vdd(vdd), .B(_1143__bF_buf6), .C(_1184_), );
  INVX2 INVX2_311 (.gnd(gnd), .A(regs_27__21_), .Y(_1185_), .vdd(vdd), );
  NAND2X1 NAND2X1_1126 (.gnd(gnd), .A(wdata[21]), .Y(_1186_), .vdd(vdd), .B(_1143__bF_buf5), );
  OAI21X1 OAI21X1_2263 (.gnd(gnd), .A(_1185_), .Y(_621_), .vdd(vdd), .B(_1143__bF_buf4), .C(_1186_), );
  INVX2 INVX2_312 (.gnd(gnd), .A(regs_27__22_), .Y(_1187_), .vdd(vdd), );
  NAND2X1 NAND2X1_1127 (.gnd(gnd), .A(wdata[22]), .Y(_1188_), .vdd(vdd), .B(_1143__bF_buf3), );
  OAI21X1 OAI21X1_2264 (.gnd(gnd), .A(_1187_), .Y(_622_), .vdd(vdd), .B(_1143__bF_buf2), .C(_1188_), );
  INVX2 INVX2_313 (.gnd(gnd), .A(regs_27__23_), .Y(_1189_), .vdd(vdd), );
  NAND2X1 NAND2X1_1128 (.gnd(gnd), .A(wdata[23]), .Y(_1190_), .vdd(vdd), .B(_1143__bF_buf1), );
  OAI21X1 OAI21X1_2265 (.gnd(gnd), .A(_1189_), .Y(_623_), .vdd(vdd), .B(_1143__bF_buf0), .C(_1190_), );
  INVX2 INVX2_314 (.gnd(gnd), .A(regs_27__24_), .Y(_1191_), .vdd(vdd), );
  NAND2X1 NAND2X1_1129 (.gnd(gnd), .A(wdata[24]), .Y(_1192_), .vdd(vdd), .B(_1143__bF_buf7), );
  OAI21X1 OAI21X1_2266 (.gnd(gnd), .A(_1191_), .Y(_624_), .vdd(vdd), .B(_1143__bF_buf6), .C(_1192_), );
  INVX2 INVX2_315 (.gnd(gnd), .A(regs_27__25_), .Y(_1193_), .vdd(vdd), );
  NAND2X1 NAND2X1_1130 (.gnd(gnd), .A(wdata[25]), .Y(_1194_), .vdd(vdd), .B(_1143__bF_buf5), );
  OAI21X1 OAI21X1_2267 (.gnd(gnd), .A(_1193_), .Y(_625_), .vdd(vdd), .B(_1143__bF_buf4), .C(_1194_), );
  INVX2 INVX2_316 (.gnd(gnd), .A(regs_27__26_), .Y(_1195_), .vdd(vdd), );
  NAND2X1 NAND2X1_1131 (.gnd(gnd), .A(wdata[26]), .Y(_1196_), .vdd(vdd), .B(_1143__bF_buf3), );
  OAI21X1 OAI21X1_2268 (.gnd(gnd), .A(_1195_), .Y(_626_), .vdd(vdd), .B(_1143__bF_buf2), .C(_1196_), );
  INVX2 INVX2_317 (.gnd(gnd), .A(regs_27__27_), .Y(_1197_), .vdd(vdd), );
  NAND2X1 NAND2X1_1132 (.gnd(gnd), .A(wdata[27]), .Y(_1198_), .vdd(vdd), .B(_1143__bF_buf1), );
  OAI21X1 OAI21X1_2269 (.gnd(gnd), .A(_1197_), .Y(_627_), .vdd(vdd), .B(_1143__bF_buf0), .C(_1198_), );
  INVX2 INVX2_318 (.gnd(gnd), .A(regs_27__28_), .Y(_1199_), .vdd(vdd), );
  NAND2X1 NAND2X1_1133 (.gnd(gnd), .A(wdata[28]), .Y(_1200_), .vdd(vdd), .B(_1143__bF_buf7), );
  OAI21X1 OAI21X1_2270 (.gnd(gnd), .A(_1199_), .Y(_628_), .vdd(vdd), .B(_1143__bF_buf6), .C(_1200_), );
  INVX2 INVX2_319 (.gnd(gnd), .A(regs_27__29_), .Y(_1201_), .vdd(vdd), );
  NAND2X1 NAND2X1_1134 (.gnd(gnd), .A(wdata[29]), .Y(_1202_), .vdd(vdd), .B(_1143__bF_buf5), );
  OAI21X1 OAI21X1_2271 (.gnd(gnd), .A(_1201_), .Y(_629_), .vdd(vdd), .B(_1143__bF_buf4), .C(_1202_), );
  INVX2 INVX2_320 (.gnd(gnd), .A(regs_27__30_), .Y(_1203_), .vdd(vdd), );
  NAND2X1 NAND2X1_1135 (.gnd(gnd), .A(wdata[30]), .Y(_1204_), .vdd(vdd), .B(_1143__bF_buf3), );
  OAI21X1 OAI21X1_2272 (.gnd(gnd), .A(_1203_), .Y(_631_), .vdd(vdd), .B(_1143__bF_buf2), .C(_1204_), );
  INVX2 INVX2_321 (.gnd(gnd), .A(regs_27__31_), .Y(_1205_), .vdd(vdd), );
  NAND2X1 NAND2X1_1136 (.gnd(gnd), .A(wdata[31]), .Y(_1206_), .vdd(vdd), .B(_1143__bF_buf1), );
  OAI21X1 OAI21X1_2273 (.gnd(gnd), .A(_1205_), .Y(_632_), .vdd(vdd), .B(_1143__bF_buf0), .C(_1206_), );
  NOR2X1 NOR2X1_285 (.gnd(gnd), .A(_1001__bF_buf9), .Y(_1207_), .vdd(vdd), .B(_1141__bF_buf2), );
  NOR2X1 NOR2X1_286 (.gnd(gnd), .A(regs_26__0_), .Y(_1208_), .vdd(vdd), .B(_1207__bF_buf7), );
  AOI21X1 AOI21X1_399 (.gnd(gnd), .A(_992__bF_buf1), .Y(_576_), .vdd(vdd), .B(_1207__bF_buf6), .C(_1208_), );
  NOR2X1 NOR2X1_287 (.gnd(gnd), .A(regs_26__1_), .Y(_1209_), .vdd(vdd), .B(_1207__bF_buf5), );
  AOI21X1 AOI21X1_400 (.gnd(gnd), .A(_1003__bF_buf1), .Y(_587_), .vdd(vdd), .B(_1207__bF_buf4), .C(_1209_), );
  NOR2X1 NOR2X1_288 (.gnd(gnd), .A(regs_26__2_), .Y(_1210_), .vdd(vdd), .B(_1207__bF_buf3), );
  AOI21X1 AOI21X1_401 (.gnd(gnd), .A(_1005__bF_buf1), .Y(_598_), .vdd(vdd), .B(_1207__bF_buf2), .C(_1210_), );
  NOR2X1 NOR2X1_289 (.gnd(gnd), .A(regs_26__3_), .Y(_1211_), .vdd(vdd), .B(_1207__bF_buf1), );
  AOI21X1 AOI21X1_402 (.gnd(gnd), .A(_1007__bF_buf1), .Y(_601_), .vdd(vdd), .B(_1207__bF_buf0), .C(_1211_), );
  NOR2X1 NOR2X1_290 (.gnd(gnd), .A(regs_26__4_), .Y(_1212_), .vdd(vdd), .B(_1207__bF_buf7), );
  AOI21X1 AOI21X1_403 (.gnd(gnd), .A(_1009__bF_buf0), .Y(_602_), .vdd(vdd), .B(_1207__bF_buf6), .C(_1212_), );
  NOR2X1 NOR2X1_291 (.gnd(gnd), .A(regs_26__5_), .Y(_1213_), .vdd(vdd), .B(_1207__bF_buf5), );
  AOI21X1 AOI21X1_404 (.gnd(gnd), .A(_1011__bF_buf0), .Y(_603_), .vdd(vdd), .B(_1207__bF_buf4), .C(_1213_), );
  NOR2X1 NOR2X1_292 (.gnd(gnd), .A(regs_26__6_), .Y(_1214_), .vdd(vdd), .B(_1207__bF_buf3), );
  AOI21X1 AOI21X1_405 (.gnd(gnd), .A(_1013__bF_buf0), .Y(_604_), .vdd(vdd), .B(_1207__bF_buf2), .C(_1214_), );
  NOR2X1 NOR2X1_293 (.gnd(gnd), .A(regs_26__7_), .Y(_1215_), .vdd(vdd), .B(_1207__bF_buf1), );
  AOI21X1 AOI21X1_406 (.gnd(gnd), .A(_1015__bF_buf0), .Y(_605_), .vdd(vdd), .B(_1207__bF_buf0), .C(_1215_), );
  NOR2X1 NOR2X1_294 (.gnd(gnd), .A(regs_26__8_), .Y(_1216_), .vdd(vdd), .B(_1207__bF_buf7), );
  AOI21X1 AOI21X1_407 (.gnd(gnd), .A(_1017__bF_buf0), .Y(_606_), .vdd(vdd), .B(_1207__bF_buf6), .C(_1216_), );
  NOR2X1 NOR2X1_295 (.gnd(gnd), .A(regs_26__9_), .Y(_1217_), .vdd(vdd), .B(_1207__bF_buf5), );
  AOI21X1 AOI21X1_408 (.gnd(gnd), .A(_1019__bF_buf0), .Y(_607_), .vdd(vdd), .B(_1207__bF_buf4), .C(_1217_), );
  NOR2X1 NOR2X1_296 (.gnd(gnd), .A(regs_26__10_), .Y(_1218_), .vdd(vdd), .B(_1207__bF_buf3), );
  AOI21X1 AOI21X1_409 (.gnd(gnd), .A(_1021__bF_buf0), .Y(_577_), .vdd(vdd), .B(_1207__bF_buf2), .C(_1218_), );
  NOR2X1 NOR2X1_297 (.gnd(gnd), .A(regs_26__11_), .Y(_1219_), .vdd(vdd), .B(_1207__bF_buf1), );
  AOI21X1 AOI21X1_410 (.gnd(gnd), .A(_1023__bF_buf0), .Y(_578_), .vdd(vdd), .B(_1207__bF_buf0), .C(_1219_), );
  NOR2X1 NOR2X1_298 (.gnd(gnd), .A(regs_26__12_), .Y(_1220_), .vdd(vdd), .B(_1207__bF_buf7), );
  AOI21X1 AOI21X1_411 (.gnd(gnd), .A(_1025__bF_buf0), .Y(_579_), .vdd(vdd), .B(_1207__bF_buf6), .C(_1220_), );
  NOR2X1 NOR2X1_299 (.gnd(gnd), .A(regs_26__13_), .Y(_1221_), .vdd(vdd), .B(_1207__bF_buf5), );
  AOI21X1 AOI21X1_412 (.gnd(gnd), .A(_1027__bF_buf0), .Y(_580_), .vdd(vdd), .B(_1207__bF_buf4), .C(_1221_), );
  NOR2X1 NOR2X1_300 (.gnd(gnd), .A(regs_26__14_), .Y(_1222_), .vdd(vdd), .B(_1207__bF_buf3), );
  AOI21X1 AOI21X1_413 (.gnd(gnd), .A(_1029__bF_buf0), .Y(_581_), .vdd(vdd), .B(_1207__bF_buf2), .C(_1222_), );
  NOR2X1 NOR2X1_301 (.gnd(gnd), .A(regs_26__15_), .Y(_1223_), .vdd(vdd), .B(_1207__bF_buf1), );
  AOI21X1 AOI21X1_414 (.gnd(gnd), .A(_1031__bF_buf0), .Y(_582_), .vdd(vdd), .B(_1207__bF_buf0), .C(_1223_), );
  NOR2X1 NOR2X1_302 (.gnd(gnd), .A(regs_26__16_), .Y(_1224_), .vdd(vdd), .B(_1207__bF_buf7), );
  AOI21X1 AOI21X1_415 (.gnd(gnd), .A(_1033__bF_buf0), .Y(_583_), .vdd(vdd), .B(_1207__bF_buf6), .C(_1224_), );
  NOR2X1 NOR2X1_303 (.gnd(gnd), .A(regs_26__17_), .Y(_1225_), .vdd(vdd), .B(_1207__bF_buf5), );
  AOI21X1 AOI21X1_416 (.gnd(gnd), .A(_1035__bF_buf0), .Y(_584_), .vdd(vdd), .B(_1207__bF_buf4), .C(_1225_), );
  NOR2X1 NOR2X1_304 (.gnd(gnd), .A(regs_26__18_), .Y(_1226_), .vdd(vdd), .B(_1207__bF_buf3), );
  AOI21X1 AOI21X1_417 (.gnd(gnd), .A(_1037__bF_buf0), .Y(_585_), .vdd(vdd), .B(_1207__bF_buf2), .C(_1226_), );
  NOR2X1 NOR2X1_305 (.gnd(gnd), .A(regs_26__19_), .Y(_1227_), .vdd(vdd), .B(_1207__bF_buf1), );
  AOI21X1 AOI21X1_418 (.gnd(gnd), .A(_1039__bF_buf0), .Y(_586_), .vdd(vdd), .B(_1207__bF_buf0), .C(_1227_), );
  NOR2X1 NOR2X1_306 (.gnd(gnd), .A(regs_26__20_), .Y(_1228_), .vdd(vdd), .B(_1207__bF_buf7), );
  AOI21X1 AOI21X1_419 (.gnd(gnd), .A(_1041__bF_buf0), .Y(_588_), .vdd(vdd), .B(_1207__bF_buf6), .C(_1228_), );
  NOR2X1 NOR2X1_307 (.gnd(gnd), .A(regs_26__21_), .Y(_1229_), .vdd(vdd), .B(_1207__bF_buf5), );
  AOI21X1 AOI21X1_420 (.gnd(gnd), .A(_1043__bF_buf0), .Y(_589_), .vdd(vdd), .B(_1207__bF_buf4), .C(_1229_), );
  NOR2X1 NOR2X1_308 (.gnd(gnd), .A(regs_26__22_), .Y(_1230_), .vdd(vdd), .B(_1207__bF_buf3), );
  AOI21X1 AOI21X1_421 (.gnd(gnd), .A(_1045__bF_buf0), .Y(_590_), .vdd(vdd), .B(_1207__bF_buf2), .C(_1230_), );
  NOR2X1 NOR2X1_309 (.gnd(gnd), .A(regs_26__23_), .Y(_1231_), .vdd(vdd), .B(_1207__bF_buf1), );
  AOI21X1 AOI21X1_422 (.gnd(gnd), .A(_1047__bF_buf0), .Y(_591_), .vdd(vdd), .B(_1207__bF_buf0), .C(_1231_), );
  NOR2X1 NOR2X1_310 (.gnd(gnd), .A(regs_26__24_), .Y(_1232_), .vdd(vdd), .B(_1207__bF_buf7), );
  AOI21X1 AOI21X1_423 (.gnd(gnd), .A(_1049__bF_buf0), .Y(_592_), .vdd(vdd), .B(_1207__bF_buf6), .C(_1232_), );
  NOR2X1 NOR2X1_311 (.gnd(gnd), .A(regs_26__25_), .Y(_1233_), .vdd(vdd), .B(_1207__bF_buf5), );
  AOI21X1 AOI21X1_424 (.gnd(gnd), .A(_1051__bF_buf0), .Y(_593_), .vdd(vdd), .B(_1207__bF_buf4), .C(_1233_), );
  NOR2X1 NOR2X1_312 (.gnd(gnd), .A(regs_26__26_), .Y(_1234_), .vdd(vdd), .B(_1207__bF_buf3), );
  AOI21X1 AOI21X1_425 (.gnd(gnd), .A(_1053__bF_buf0), .Y(_594_), .vdd(vdd), .B(_1207__bF_buf2), .C(_1234_), );
  NOR2X1 NOR2X1_313 (.gnd(gnd), .A(regs_26__27_), .Y(_1235_), .vdd(vdd), .B(_1207__bF_buf1), );
  AOI21X1 AOI21X1_426 (.gnd(gnd), .A(_1055__bF_buf0), .Y(_595_), .vdd(vdd), .B(_1207__bF_buf0), .C(_1235_), );
  NOR2X1 NOR2X1_314 (.gnd(gnd), .A(regs_26__28_), .Y(_1236_), .vdd(vdd), .B(_1207__bF_buf7), );
  AOI21X1 AOI21X1_427 (.gnd(gnd), .A(_1057__bF_buf0), .Y(_596_), .vdd(vdd), .B(_1207__bF_buf6), .C(_1236_), );
  NOR2X1 NOR2X1_315 (.gnd(gnd), .A(regs_26__29_), .Y(_1237_), .vdd(vdd), .B(_1207__bF_buf5), );
  AOI21X1 AOI21X1_428 (.gnd(gnd), .A(_1059__bF_buf0), .Y(_597_), .vdd(vdd), .B(_1207__bF_buf4), .C(_1237_), );
  NOR2X1 NOR2X1_316 (.gnd(gnd), .A(regs_26__30_), .Y(_1238_), .vdd(vdd), .B(_1207__bF_buf3), );
  AOI21X1 AOI21X1_429 (.gnd(gnd), .A(_1061__bF_buf0), .Y(_599_), .vdd(vdd), .B(_1207__bF_buf2), .C(_1238_), );
  NOR2X1 NOR2X1_317 (.gnd(gnd), .A(regs_26__31_), .Y(_1239_), .vdd(vdd), .B(_1207__bF_buf1), );
  AOI21X1 AOI21X1_430 (.gnd(gnd), .A(_1063__bF_buf0), .Y(_600_), .vdd(vdd), .B(_1207__bF_buf0), .C(_1239_), );
  NAND2X1 NAND2X1_1137 (.gnd(gnd), .A(_1068_), .Y(_1240_), .vdd(vdd), .B(_1140_), );
  OAI21X1 OAI21X1_2274 (.gnd(gnd), .A(_1141__bF_buf1), .Y(_1241_), .vdd(vdd), .B(_1070__bF_buf9), .C(regs_25__0_), );
  OAI21X1 OAI21X1_2275 (.gnd(gnd), .A(_992__bF_buf0), .Y(_544_), .vdd(vdd), .B(_1240__bF_buf4), .C(_1241_), );
  OAI21X1 OAI21X1_2276 (.gnd(gnd), .A(_1141__bF_buf0), .Y(_1242_), .vdd(vdd), .B(_1070__bF_buf8), .C(regs_25__1_), );
  OAI21X1 OAI21X1_2277 (.gnd(gnd), .A(_1003__bF_buf0), .Y(_555_), .vdd(vdd), .B(_1240__bF_buf3), .C(_1242_), );
  OAI21X1 OAI21X1_2278 (.gnd(gnd), .A(_1141__bF_buf7), .Y(_1243_), .vdd(vdd), .B(_1070__bF_buf7), .C(regs_25__2_), );
  OAI21X1 OAI21X1_2279 (.gnd(gnd), .A(_1005__bF_buf0), .Y(_566_), .vdd(vdd), .B(_1240__bF_buf2), .C(_1243_), );
  OAI21X1 OAI21X1_2280 (.gnd(gnd), .A(_1141__bF_buf6), .Y(_1244_), .vdd(vdd), .B(_1070__bF_buf6), .C(regs_25__3_), );
  OAI21X1 OAI21X1_2281 (.gnd(gnd), .A(_1007__bF_buf0), .Y(_569_), .vdd(vdd), .B(_1240__bF_buf1), .C(_1244_), );
  OAI21X1 OAI21X1_2282 (.gnd(gnd), .A(_1141__bF_buf5), .Y(_1245_), .vdd(vdd), .B(_1070__bF_buf5), .C(regs_25__4_), );
  OAI21X1 OAI21X1_2283 (.gnd(gnd), .A(_1009__bF_buf3), .Y(_570_), .vdd(vdd), .B(_1240__bF_buf0), .C(_1245_), );
  OAI21X1 OAI21X1_2284 (.gnd(gnd), .A(_1141__bF_buf4), .Y(_1246_), .vdd(vdd), .B(_1070__bF_buf4), .C(regs_25__5_), );
  OAI21X1 OAI21X1_2285 (.gnd(gnd), .A(_1011__bF_buf3), .Y(_571_), .vdd(vdd), .B(_1240__bF_buf4), .C(_1246_), );
  OAI21X1 OAI21X1_2286 (.gnd(gnd), .A(_1141__bF_buf3), .Y(_1247_), .vdd(vdd), .B(_1070__bF_buf3), .C(regs_25__6_), );
  OAI21X1 OAI21X1_2287 (.gnd(gnd), .A(_1013__bF_buf3), .Y(_572_), .vdd(vdd), .B(_1240__bF_buf3), .C(_1247_), );
  OAI21X1 OAI21X1_2288 (.gnd(gnd), .A(_1141__bF_buf2), .Y(_1248_), .vdd(vdd), .B(_1070__bF_buf2), .C(regs_25__7_), );
  OAI21X1 OAI21X1_2289 (.gnd(gnd), .A(_1015__bF_buf3), .Y(_573_), .vdd(vdd), .B(_1240__bF_buf2), .C(_1248_), );
  OAI21X1 OAI21X1_2290 (.gnd(gnd), .A(_1141__bF_buf1), .Y(_1249_), .vdd(vdd), .B(_1070__bF_buf1), .C(regs_25__8_), );
  OAI21X1 OAI21X1_2291 (.gnd(gnd), .A(_1017__bF_buf3), .Y(_574_), .vdd(vdd), .B(_1240__bF_buf1), .C(_1249_), );
  OAI21X1 OAI21X1_2292 (.gnd(gnd), .A(_1141__bF_buf0), .Y(_1250_), .vdd(vdd), .B(_1070__bF_buf0), .C(regs_25__9_), );
  OAI21X1 OAI21X1_2293 (.gnd(gnd), .A(_1019__bF_buf3), .Y(_575_), .vdd(vdd), .B(_1240__bF_buf0), .C(_1250_), );
  OAI21X1 OAI21X1_2294 (.gnd(gnd), .A(_1141__bF_buf7), .Y(_1251_), .vdd(vdd), .B(_1070__bF_buf10), .C(regs_25__10_), );
  OAI21X1 OAI21X1_2295 (.gnd(gnd), .A(_1021__bF_buf3), .Y(_545_), .vdd(vdd), .B(_1240__bF_buf4), .C(_1251_), );
  OAI21X1 OAI21X1_2296 (.gnd(gnd), .A(_1141__bF_buf6), .Y(_1252_), .vdd(vdd), .B(_1070__bF_buf9), .C(regs_25__11_), );
  OAI21X1 OAI21X1_2297 (.gnd(gnd), .A(_1023__bF_buf3), .Y(_546_), .vdd(vdd), .B(_1240__bF_buf3), .C(_1252_), );
  OAI21X1 OAI21X1_2298 (.gnd(gnd), .A(_1141__bF_buf5), .Y(_1253_), .vdd(vdd), .B(_1070__bF_buf8), .C(regs_25__12_), );
  OAI21X1 OAI21X1_2299 (.gnd(gnd), .A(_1025__bF_buf3), .Y(_547_), .vdd(vdd), .B(_1240__bF_buf2), .C(_1253_), );
  OAI21X1 OAI21X1_2300 (.gnd(gnd), .A(_1141__bF_buf4), .Y(_1254_), .vdd(vdd), .B(_1070__bF_buf7), .C(regs_25__13_), );
  OAI21X1 OAI21X1_2301 (.gnd(gnd), .A(_1027__bF_buf3), .Y(_548_), .vdd(vdd), .B(_1240__bF_buf1), .C(_1254_), );
  OAI21X1 OAI21X1_2302 (.gnd(gnd), .A(_1141__bF_buf3), .Y(_1255_), .vdd(vdd), .B(_1070__bF_buf6), .C(regs_25__14_), );
  OAI21X1 OAI21X1_2303 (.gnd(gnd), .A(_1029__bF_buf3), .Y(_549_), .vdd(vdd), .B(_1240__bF_buf0), .C(_1255_), );
  OAI21X1 OAI21X1_2304 (.gnd(gnd), .A(_1141__bF_buf2), .Y(_1256_), .vdd(vdd), .B(_1070__bF_buf5), .C(regs_25__15_), );
  OAI21X1 OAI21X1_2305 (.gnd(gnd), .A(_1031__bF_buf3), .Y(_550_), .vdd(vdd), .B(_1240__bF_buf4), .C(_1256_), );
  OAI21X1 OAI21X1_2306 (.gnd(gnd), .A(_1141__bF_buf1), .Y(_1257_), .vdd(vdd), .B(_1070__bF_buf4), .C(regs_25__16_), );
  OAI21X1 OAI21X1_2307 (.gnd(gnd), .A(_1033__bF_buf3), .Y(_551_), .vdd(vdd), .B(_1240__bF_buf3), .C(_1257_), );
  OAI21X1 OAI21X1_2308 (.gnd(gnd), .A(_1141__bF_buf0), .Y(_1258_), .vdd(vdd), .B(_1070__bF_buf3), .C(regs_25__17_), );
  OAI21X1 OAI21X1_2309 (.gnd(gnd), .A(_1035__bF_buf3), .Y(_552_), .vdd(vdd), .B(_1240__bF_buf2), .C(_1258_), );
  OAI21X1 OAI21X1_2310 (.gnd(gnd), .A(_1141__bF_buf7), .Y(_1259_), .vdd(vdd), .B(_1070__bF_buf2), .C(regs_25__18_), );
  OAI21X1 OAI21X1_2311 (.gnd(gnd), .A(_1037__bF_buf3), .Y(_553_), .vdd(vdd), .B(_1240__bF_buf1), .C(_1259_), );
  OAI21X1 OAI21X1_2312 (.gnd(gnd), .A(_1141__bF_buf6), .Y(_1260_), .vdd(vdd), .B(_1070__bF_buf1), .C(regs_25__19_), );
  OAI21X1 OAI21X1_2313 (.gnd(gnd), .A(_1039__bF_buf3), .Y(_554_), .vdd(vdd), .B(_1240__bF_buf0), .C(_1260_), );
  OAI21X1 OAI21X1_2314 (.gnd(gnd), .A(_1141__bF_buf5), .Y(_1261_), .vdd(vdd), .B(_1070__bF_buf0), .C(regs_25__20_), );
  OAI21X1 OAI21X1_2315 (.gnd(gnd), .A(_1041__bF_buf3), .Y(_556_), .vdd(vdd), .B(_1240__bF_buf4), .C(_1261_), );
  OAI21X1 OAI21X1_2316 (.gnd(gnd), .A(_1141__bF_buf4), .Y(_1262_), .vdd(vdd), .B(_1070__bF_buf10), .C(regs_25__21_), );
  OAI21X1 OAI21X1_2317 (.gnd(gnd), .A(_1043__bF_buf3), .Y(_557_), .vdd(vdd), .B(_1240__bF_buf3), .C(_1262_), );
  OAI21X1 OAI21X1_2318 (.gnd(gnd), .A(_1141__bF_buf3), .Y(_1263_), .vdd(vdd), .B(_1070__bF_buf9), .C(regs_25__22_), );
  OAI21X1 OAI21X1_2319 (.gnd(gnd), .A(_1045__bF_buf3), .Y(_558_), .vdd(vdd), .B(_1240__bF_buf2), .C(_1263_), );
  OAI21X1 OAI21X1_2320 (.gnd(gnd), .A(_1141__bF_buf2), .Y(_1264_), .vdd(vdd), .B(_1070__bF_buf8), .C(regs_25__23_), );
  OAI21X1 OAI21X1_2321 (.gnd(gnd), .A(_1047__bF_buf3), .Y(_559_), .vdd(vdd), .B(_1240__bF_buf1), .C(_1264_), );
  OAI21X1 OAI21X1_2322 (.gnd(gnd), .A(_1141__bF_buf1), .Y(_1265_), .vdd(vdd), .B(_1070__bF_buf7), .C(regs_25__24_), );
  OAI21X1 OAI21X1_2323 (.gnd(gnd), .A(_1049__bF_buf3), .Y(_560_), .vdd(vdd), .B(_1240__bF_buf0), .C(_1265_), );
  OAI21X1 OAI21X1_2324 (.gnd(gnd), .A(_1141__bF_buf0), .Y(_1266_), .vdd(vdd), .B(_1070__bF_buf6), .C(regs_25__25_), );
  OAI21X1 OAI21X1_2325 (.gnd(gnd), .A(_1051__bF_buf3), .Y(_561_), .vdd(vdd), .B(_1240__bF_buf4), .C(_1266_), );
  OAI21X1 OAI21X1_2326 (.gnd(gnd), .A(_1141__bF_buf7), .Y(_1267_), .vdd(vdd), .B(_1070__bF_buf5), .C(regs_25__26_), );
  OAI21X1 OAI21X1_2327 (.gnd(gnd), .A(_1053__bF_buf3), .Y(_562_), .vdd(vdd), .B(_1240__bF_buf3), .C(_1267_), );
  OAI21X1 OAI21X1_2328 (.gnd(gnd), .A(_1141__bF_buf6), .Y(_1268_), .vdd(vdd), .B(_1070__bF_buf4), .C(regs_25__27_), );
  OAI21X1 OAI21X1_2329 (.gnd(gnd), .A(_1055__bF_buf3), .Y(_563_), .vdd(vdd), .B(_1240__bF_buf2), .C(_1268_), );
  OAI21X1 OAI21X1_2330 (.gnd(gnd), .A(_1141__bF_buf5), .Y(_1269_), .vdd(vdd), .B(_1070__bF_buf3), .C(regs_25__28_), );
  OAI21X1 OAI21X1_2331 (.gnd(gnd), .A(_1057__bF_buf3), .Y(_564_), .vdd(vdd), .B(_1240__bF_buf1), .C(_1269_), );
  OAI21X1 OAI21X1_2332 (.gnd(gnd), .A(_1141__bF_buf4), .Y(_1270_), .vdd(vdd), .B(_1070__bF_buf2), .C(regs_25__29_), );
  OAI21X1 OAI21X1_2333 (.gnd(gnd), .A(_1059__bF_buf3), .Y(_565_), .vdd(vdd), .B(_1240__bF_buf0), .C(_1270_), );
  OAI21X1 OAI21X1_2334 (.gnd(gnd), .A(_1141__bF_buf3), .Y(_1271_), .vdd(vdd), .B(_1070__bF_buf1), .C(regs_25__30_), );
  OAI21X1 OAI21X1_2335 (.gnd(gnd), .A(_1061__bF_buf3), .Y(_567_), .vdd(vdd), .B(_1240__bF_buf4), .C(_1271_), );
  OAI21X1 OAI21X1_2336 (.gnd(gnd), .A(_1141__bF_buf2), .Y(_1272_), .vdd(vdd), .B(_1070__bF_buf0), .C(regs_25__31_), );
  OAI21X1 OAI21X1_2337 (.gnd(gnd), .A(_1063__bF_buf3), .Y(_568_), .vdd(vdd), .B(_1240__bF_buf3), .C(_1272_), );
  INVX1 INVX1_167 (.gnd(gnd), .A(_1104__bF_buf14), .Y(_1273_), .vdd(vdd), );
  NAND2X1 NAND2X1_1138 (.gnd(gnd), .A(_1140_), .Y(_1274_), .vdd(vdd), .B(_1273_), );
  OAI21X1 OAI21X1_2338 (.gnd(gnd), .A(_1141__bF_buf1), .Y(_1275_), .vdd(vdd), .B(_1104__bF_buf13), .C(regs_24__0_), );
  OAI21X1 OAI21X1_2339 (.gnd(gnd), .A(_1274__bF_buf1), .Y(_512_), .vdd(vdd), .B(_992__bF_buf3), .C(_1275_), );
  OAI21X1 OAI21X1_2340 (.gnd(gnd), .A(_1141__bF_buf0), .Y(_1276_), .vdd(vdd), .B(_1104__bF_buf12), .C(regs_24__1_), );
  OAI21X1 OAI21X1_2341 (.gnd(gnd), .A(_1274__bF_buf0), .Y(_523_), .vdd(vdd), .B(_1003__bF_buf3), .C(_1276_), );
  OAI21X1 OAI21X1_2342 (.gnd(gnd), .A(_1141__bF_buf7), .Y(_1277_), .vdd(vdd), .B(_1104__bF_buf11), .C(regs_24__2_), );
  OAI21X1 OAI21X1_2343 (.gnd(gnd), .A(_1274__bF_buf4), .Y(_534_), .vdd(vdd), .B(_1005__bF_buf3), .C(_1277_), );
  OAI21X1 OAI21X1_2344 (.gnd(gnd), .A(_1141__bF_buf6), .Y(_1278_), .vdd(vdd), .B(_1104__bF_buf10), .C(regs_24__3_), );
  OAI21X1 OAI21X1_2345 (.gnd(gnd), .A(_1274__bF_buf3), .Y(_537_), .vdd(vdd), .B(_1007__bF_buf3), .C(_1278_), );
  CLKBUF3 CLKBUF3__1 (.A(clk_bF_buf89), .Y(random_clk_bf3__1), );
  CLKBUF3 CLKBUF3__2 (.Y(random_clk_bf3__2), .A(clk_bF_buf89), );
  CLKBUF3 CLKBUF3__21 (.A(clk_bF_buf80), .Y(random_clk_bf3__21), );
  CLKBUF3 CLKBUF3__22 (.Y(random_clk_bf3__22), .A(clk_bF_buf80), );
  CLKBUF3 CLKBUF3__41 (.A(clk_bF_buf71), .Y(random_clk_bf3__41), );
  CLKBUF3 CLKBUF3__42 (.Y(random_clk_bf3__42), .A(clk_bF_buf71), );
  CLKBUF3 CLKBUF3__61 (.A(clk_bF_buf62), .Y(random_clk_bf3__61), );
  CLKBUF3 CLKBUF3__62 (.Y(random_clk_bf3__62), .A(clk_bF_buf62), );
  CLKBUF3 CLKBUF3__81 (.A(clk_bF_buf53), .Y(random_clk_bf3__81), );
  CLKBUF3 CLKBUF3__82 (.Y(random_clk_bf3__82), .A(clk_bF_buf53), );
  CLKBUF3 CLKBUF3__101 (.A(clk_bF_buf44), .Y(random_clk_bf3__101), );
  CLKBUF3 CLKBUF3__102 (.Y(random_clk_bf3__102), .A(clk_bF_buf44), );
  CLKBUF3 CLKBUF3__121 (.A(clk_bF_buf35), .Y(random_clk_bf3__121), );
  CLKBUF3 CLKBUF3__122 (.Y(random_clk_bf3__122), .A(clk_bF_buf35), );
  CLKBUF3 CLKBUF3__141 (.A(clk_bF_buf26), .Y(random_clk_bf3__141), );
  CLKBUF3 CLKBUF3__142 (.Y(random_clk_bf3__142), .A(clk_bF_buf26), );
  CLKBUF3 CLKBUF3__161 (.A(clk_bF_buf17), .Y(random_clk_bf3__161), );
  CLKBUF3 CLKBUF3__162 (.Y(random_clk_bf3__162), .A(clk_bF_buf17), );
  CLKBUF3 CLKBUF3__181 (.A(clk_bF_buf8), .Y(random_clk_bf3__181), );
  CLKBUF3 CLKBUF3__182 (.Y(random_clk_bf3__182), .A(clk_bF_buf8), );
  CLKBUF3 CLKBUF3__201 (.A(clk_bF_buf88), .Y(random_clk_bf3__201), );
  CLKBUF3 CLKBUF3__202 (.Y(random_clk_bf3__202), .A(clk_bF_buf88), );
  CLKBUF3 CLKBUF3__221 (.A(clk_bF_buf79), .Y(random_clk_bf3__221), );
  CLKBUF3 CLKBUF3__222 (.Y(random_clk_bf3__222), .A(clk_bF_buf79), );
  CLKBUF3 CLKBUF3__241 (.A(clk_bF_buf70), .Y(random_clk_bf3__241), );
  CLKBUF3 CLKBUF3__242 (.Y(random_clk_bf3__242), .A(clk_bF_buf70), );
  CLKBUF3 CLKBUF3__261 (.A(clk_bF_buf61), .Y(random_clk_bf3__261), );
  CLKBUF3 CLKBUF3__262 (.Y(random_clk_bf3__262), .A(clk_bF_buf61), );
  CLKBUF3 CLKBUF3__281 (.A(clk_bF_buf52), .Y(random_clk_bf3__281), );
  CLKBUF3 CLKBUF3__282 (.Y(random_clk_bf3__282), .A(clk_bF_buf52), );
  CLKBUF3 CLKBUF3__301 (.A(clk_bF_buf43), .Y(random_clk_bf3__301), );
  CLKBUF3 CLKBUF3__302 (.Y(random_clk_bf3__302), .A(clk_bF_buf43), );
  CLKBUF3 CLKBUF3__321 (.A(clk_bF_buf34), .Y(random_clk_bf3__321), );
  CLKBUF3 CLKBUF3__322 (.Y(random_clk_bf3__322), .A(clk_bF_buf34), );
  CLKBUF3 CLKBUF3__341 (.A(clk_bF_buf25), .Y(random_clk_bf3__341), );
  CLKBUF3 CLKBUF3__342 (.Y(random_clk_bf3__342), .A(clk_bF_buf25), );
  CLKBUF3 CLKBUF3__361 (.A(clk_bF_buf16), .Y(random_clk_bf3__361), );
  CLKBUF3 CLKBUF3__362 (.Y(random_clk_bf3__362), .A(clk_bF_buf16), );
  CLKBUF3 CLKBUF3__381 (.A(clk_bF_buf7), .Y(random_clk_bf3__381), );
  CLKBUF3 CLKBUF3__382 (.Y(random_clk_bf3__382), .A(clk_bF_buf7), );
  CLKBUF3 CLKBUF3__401 (.A(clk_bF_buf96), .Y(random_clk_bf3__401), );
  CLKBUF3 CLKBUF3__402 (.Y(random_clk_bf3__402), .A(clk_bF_buf96), );
  CLKBUF3 CLKBUF3__421 (.A(clk_bF_buf87), .Y(random_clk_bf3__421), );
  CLKBUF3 CLKBUF3__422 (.Y(random_clk_bf3__422), .A(clk_bF_buf87), );
  CLKBUF3 CLKBUF3__441 (.A(clk_bF_buf78), .Y(random_clk_bf3__441), );
  CLKBUF3 CLKBUF3__442 (.Y(random_clk_bf3__442), .A(clk_bF_buf78), );
  CLKBUF3 CLKBUF3__461 (.A(clk_bF_buf69), .Y(random_clk_bf3__461), );
  CLKBUF3 CLKBUF3__462 (.Y(random_clk_bf3__462), .A(clk_bF_buf69), );
  CLKBUF3 CLKBUF3__481 (.A(clk_bF_buf60), .Y(random_clk_bf3__481), );
  CLKBUF3 CLKBUF3__482 (.Y(random_clk_bf3__482), .A(clk_bF_buf60), );
  CLKBUF3 CLKBUF3__501 (.A(clk_bF_buf51), .Y(random_clk_bf3__501), );
  CLKBUF3 CLKBUF3__502 (.Y(random_clk_bf3__502), .A(clk_bF_buf51), );
  CLKBUF3 CLKBUF3__521 (.A(clk_bF_buf42), .Y(random_clk_bf3__521), );
  CLKBUF3 CLKBUF3__522 (.Y(random_clk_bf3__522), .A(clk_bF_buf42), );
  CLKBUF3 CLKBUF3__541 (.A(clk_bF_buf33), .Y(random_clk_bf3__541), );
  CLKBUF3 CLKBUF3__542 (.Y(random_clk_bf3__542), .A(clk_bF_buf33), );
  CLKBUF3 CLKBUF3__561 (.A(clk_bF_buf24), .Y(random_clk_bf3__561), );
  CLKBUF3 CLKBUF3__562 (.Y(random_clk_bf3__562), .A(clk_bF_buf24), );
  CLKBUF3 CLKBUF3__581 (.A(clk_bF_buf15), .Y(random_clk_bf3__581), );
  CLKBUF3 CLKBUF3__582 (.Y(random_clk_bf3__582), .A(clk_bF_buf15), );
  CLKBUF3 CLKBUF3__601 (.A(clk_bF_buf6), .Y(random_clk_bf3__601), );
  CLKBUF3 CLKBUF3__602 (.Y(random_clk_bf3__602), .A(clk_bF_buf6), );
  CLKBUF3 CLKBUF3__621 (.A(clk_bF_buf95), .Y(random_clk_bf3__621), );
  CLKBUF3 CLKBUF3__622 (.Y(random_clk_bf3__622), .A(clk_bF_buf95), );
  CLKBUF3 CLKBUF3__641 (.A(clk_bF_buf86), .Y(random_clk_bf3__641), );
  CLKBUF3 CLKBUF3__642 (.Y(random_clk_bf3__642), .A(clk_bF_buf86), );
  CLKBUF3 CLKBUF3__661 (.A(clk_bF_buf77), .Y(random_clk_bf3__661), );
  CLKBUF3 CLKBUF3__662 (.Y(random_clk_bf3__662), .A(clk_bF_buf77), );
  CLKBUF3 CLKBUF3__681 (.A(clk_bF_buf68), .Y(random_clk_bf3__681), );
  CLKBUF3 CLKBUF3__682 (.Y(random_clk_bf3__682), .A(clk_bF_buf68), );
  CLKBUF3 CLKBUF3__701 (.A(clk_bF_buf59), .Y(random_clk_bf3__701), );
  CLKBUF3 CLKBUF3__702 (.Y(random_clk_bf3__702), .A(clk_bF_buf59), );
  CLKBUF3 CLKBUF3__721 (.A(clk_bF_buf50), .Y(random_clk_bf3__721), );
  CLKBUF3 CLKBUF3__722 (.Y(random_clk_bf3__722), .A(clk_bF_buf50), );
  CLKBUF3 CLKBUF3__741 (.A(clk_bF_buf41), .Y(random_clk_bf3__741), );
  CLKBUF3 CLKBUF3__742 (.Y(random_clk_bf3__742), .A(clk_bF_buf41), );
  CLKBUF3 CLKBUF3__761 (.A(clk_bF_buf32), .Y(random_clk_bf3__761), );
  CLKBUF3 CLKBUF3__762 (.Y(random_clk_bf3__762), .A(clk_bF_buf32), );
  CLKBUF3 CLKBUF3__781 (.A(clk_bF_buf23), .Y(random_clk_bf3__781), );
  CLKBUF3 CLKBUF3__782 (.Y(random_clk_bf3__782), .A(clk_bF_buf23), );
  CLKBUF3 CLKBUF3__801 (.A(clk_bF_buf14), .Y(random_clk_bf3__801), );
  CLKBUF3 CLKBUF3__802 (.Y(random_clk_bf3__802), .A(clk_bF_buf14), );
  CLKBUF3 CLKBUF3__821 (.A(clk_bF_buf5), .Y(random_clk_bf3__821), );
  CLKBUF3 CLKBUF3__822 (.Y(random_clk_bf3__822), .A(clk_bF_buf5), );
  CLKBUF3 CLKBUF3__841 (.A(clk_bF_buf94), .Y(random_clk_bf3__841), );
  CLKBUF3 CLKBUF3__842 (.Y(random_clk_bf3__842), .A(clk_bF_buf94), );
  CLKBUF3 CLKBUF3__861 (.A(clk_bF_buf85), .Y(random_clk_bf3__861), );
  CLKBUF3 CLKBUF3__862 (.Y(random_clk_bf3__862), .A(clk_bF_buf85), );
  CLKBUF3 CLKBUF3__881 (.A(clk_bF_buf76), .Y(random_clk_bf3__881), );
  CLKBUF3 CLKBUF3__882 (.Y(random_clk_bf3__882), .A(clk_bF_buf76), );
  CLKBUF3 CLKBUF3__901 (.A(clk_bF_buf67), .Y(random_clk_bf3__901), );
  CLKBUF3 CLKBUF3__902 (.Y(random_clk_bf3__902), .A(clk_bF_buf67), );
  CLKBUF3 CLKBUF3__921 (.A(clk_bF_buf58), .Y(random_clk_bf3__921), );
  CLKBUF3 CLKBUF3__922 (.Y(random_clk_bf3__922), .A(clk_bF_buf58), );
  CLKBUF3 CLKBUF3__941 (.A(clk_bF_buf49), .Y(random_clk_bf3__941), );
  CLKBUF3 CLKBUF3__942 (.Y(random_clk_bf3__942), .A(clk_bF_buf49), );
  CLKBUF3 CLKBUF3__961 (.A(clk_bF_buf40), .Y(random_clk_bf3__961), );
  CLKBUF3 CLKBUF3__962 (.Y(random_clk_bf3__962), .A(clk_bF_buf40), );
  CLKBUF3 CLKBUF3__981 (.A(clk_bF_buf31), .Y(random_clk_bf3__981), );
  CLKBUF3 CLKBUF3__982 (.Y(random_clk_bf3__982), .A(clk_bF_buf31), );
  CLKBUF3 CLKBUF3__1001 (.A(clk_bF_buf22), .Y(random_clk_bf3__1001), );
  CLKBUF3 CLKBUF3__1002 (.Y(random_clk_bf3__1002), .A(clk_bF_buf22), );
  CLKBUF3 CLKBUF3__1021 (.A(clk_bF_buf13), .Y(random_clk_bf3__1021), );
  CLKBUF3 CLKBUF3__1022 (.Y(random_clk_bf3__1022), .A(clk_bF_buf13), );
  CLKBUF3 CLKBUF3__1041 (.A(clk_bF_buf4), .Y(random_clk_bf3__1041), );
  CLKBUF3 CLKBUF3__1042 (.Y(random_clk_bf3__1042), .A(clk_bF_buf4), );
  CLKBUF3 CLKBUF3__1061 (.A(clk_bF_buf93), .Y(random_clk_bf3__1061), );
  CLKBUF3 CLKBUF3__1062 (.Y(random_clk_bf3__1062), .A(clk_bF_buf93), );
  CLKBUF3 CLKBUF3__1081 (.A(clk_bF_buf84), .Y(random_clk_bf3__1081), );
  CLKBUF3 CLKBUF3__1082 (.Y(random_clk_bf3__1082), .A(clk_bF_buf84), );
  CLKBUF3 CLKBUF3__1101 (.A(clk_bF_buf75), .Y(random_clk_bf3__1101), );
  CLKBUF3 CLKBUF3__1102 (.Y(random_clk_bf3__1102), .A(clk_bF_buf75), );
  CLKBUF3 CLKBUF3__1121 (.A(clk_bF_buf66), .Y(random_clk_bf3__1121), );
  CLKBUF3 CLKBUF3__1122 (.Y(random_clk_bf3__1122), .A(clk_bF_buf66), );
  CLKBUF3 CLKBUF3__1141 (.A(clk_bF_buf57), .Y(random_clk_bf3__1141), );
  CLKBUF3 CLKBUF3__1142 (.Y(random_clk_bf3__1142), .A(clk_bF_buf57), );
  CLKBUF3 CLKBUF3__1161 (.A(clk_bF_buf48), .Y(random_clk_bf3__1161), );
  CLKBUF3 CLKBUF3__1162 (.Y(random_clk_bf3__1162), .A(clk_bF_buf48), );
  CLKBUF3 CLKBUF3__1181 (.A(clk_bF_buf39), .Y(random_clk_bf3__1181), );
  CLKBUF3 CLKBUF3__1182 (.Y(random_clk_bf3__1182), .A(clk_bF_buf39), );
  CLKBUF3 CLKBUF3__1201 (.A(clk_bF_buf30), .Y(random_clk_bf3__1201), );
  CLKBUF3 CLKBUF3__1202 (.Y(random_clk_bf3__1202), .A(clk_bF_buf30), );
  CLKBUF3 CLKBUF3__1221 (.A(clk_bF_buf21), .Y(random_clk_bf3__1221), );
  CLKBUF3 CLKBUF3__1222 (.Y(random_clk_bf3__1222), .A(clk_bF_buf21), );
  CLKBUF3 CLKBUF3__1241 (.A(clk_bF_buf12), .Y(random_clk_bf3__1241), );
  CLKBUF3 CLKBUF3__1242 (.Y(random_clk_bf3__1242), .A(clk_bF_buf12), );
  CLKBUF3 CLKBUF3__1261 (.A(clk_bF_buf3), .Y(random_clk_bf3__1261), );
  CLKBUF3 CLKBUF3__1262 (.Y(random_clk_bf3__1262), .A(clk_bF_buf3), );
  CLKBUF3 CLKBUF3__1281 (.A(clk_bF_buf92), .Y(random_clk_bf3__1281), );
  CLKBUF3 CLKBUF3__1282 (.Y(random_clk_bf3__1282), .A(clk_bF_buf92), );
  CLKBUF3 CLKBUF3__1301 (.A(clk_bF_buf83), .Y(random_clk_bf3__1301), );
  CLKBUF3 CLKBUF3__1302 (.Y(random_clk_bf3__1302), .A(clk_bF_buf83), );
  CLKBUF3 CLKBUF3__1321 (.A(clk_bF_buf74), .Y(random_clk_bf3__1321), );
  CLKBUF3 CLKBUF3__1322 (.Y(random_clk_bf3__1322), .A(clk_bF_buf74), );
  CLKBUF3 CLKBUF3__1341 (.A(clk_bF_buf65), .Y(random_clk_bf3__1341), );
  CLKBUF3 CLKBUF3__1342 (.Y(random_clk_bf3__1342), .A(clk_bF_buf65), );
  CLKBUF3 CLKBUF3__1361 (.A(clk_bF_buf56), .Y(random_clk_bf3__1361), );
  CLKBUF3 CLKBUF3__1362 (.Y(random_clk_bf3__1362), .A(clk_bF_buf56), );
  CLKBUF3 CLKBUF3__1381 (.A(clk_bF_buf47), .Y(random_clk_bf3__1381), );
  CLKBUF3 CLKBUF3__1382 (.Y(random_clk_bf3__1382), .A(clk_bF_buf47), );
  CLKBUF3 CLKBUF3__1401 (.A(clk_bF_buf38), .Y(random_clk_bf3__1401), );
  CLKBUF3 CLKBUF3__1402 (.Y(random_clk_bf3__1402), .A(clk_bF_buf38), );
  CLKBUF3 CLKBUF3__1421 (.A(clk_bF_buf29), .Y(random_clk_bf3__1421), );
  CLKBUF3 CLKBUF3__1422 (.Y(random_clk_bf3__1422), .A(clk_bF_buf29), );
  CLKBUF3 CLKBUF3__1441 (.A(clk_bF_buf20), .Y(random_clk_bf3__1441), );
  CLKBUF3 CLKBUF3__1442 (.Y(random_clk_bf3__1442), .A(clk_bF_buf20), );
  CLKBUF3 CLKBUF3__1461 (.A(clk_bF_buf11), .Y(random_clk_bf3__1461), );
  CLKBUF3 CLKBUF3__1462 (.Y(random_clk_bf3__1462), .A(clk_bF_buf11), );
  CLKBUF3 CLKBUF3__1481 (.A(clk_bF_buf2), .Y(random_clk_bf3__1481), );
  CLKBUF3 CLKBUF3__1482 (.Y(random_clk_bf3__1482), .A(clk_bF_buf2), );
  CLKBUF3 CLKBUF3__1501 (.A(clk_bF_buf91), .Y(random_clk_bf3__1501), );
  CLKBUF3 CLKBUF3__1502 (.Y(random_clk_bf3__1502), .A(clk_bF_buf91), );
  CLKBUF3 CLKBUF3__1521 (.A(clk_bF_buf82), .Y(random_clk_bf3__1521), );
  CLKBUF3 CLKBUF3__1522 (.Y(random_clk_bf3__1522), .A(clk_bF_buf82), );
  CLKBUF3 CLKBUF3__1541 (.A(clk_bF_buf73), .Y(random_clk_bf3__1541), );
  CLKBUF3 CLKBUF3__1542 (.Y(random_clk_bf3__1542), .A(clk_bF_buf73), );
  CLKBUF3 CLKBUF3__1561 (.A(clk_bF_buf64), .Y(random_clk_bf3__1561), );
  CLKBUF3 CLKBUF3__1562 (.Y(random_clk_bf3__1562), .A(clk_bF_buf64), );
  CLKBUF3 CLKBUF3__1581 (.A(clk_bF_buf55), .Y(random_clk_bf3__1581), );
  CLKBUF3 CLKBUF3__1582 (.Y(random_clk_bf3__1582), .A(clk_bF_buf55), );
  CLKBUF3 CLKBUF3__1601 (.A(clk_bF_buf46), .Y(random_clk_bf3__1601), );
  CLKBUF3 CLKBUF3__1602 (.Y(random_clk_bf3__1602), .A(clk_bF_buf46), );
  CLKBUF3 CLKBUF3__1621 (.A(clk_bF_buf37), .Y(random_clk_bf3__1621), );
  CLKBUF3 CLKBUF3__1622 (.Y(random_clk_bf3__1622), .A(clk_bF_buf37), );
  CLKBUF3 CLKBUF3__1641 (.A(clk_bF_buf28), .Y(random_clk_bf3__1641), );
  CLKBUF3 CLKBUF3__1642 (.Y(random_clk_bf3__1642), .A(clk_bF_buf28), );
  CLKBUF3 CLKBUF3__1661 (.A(clk_bF_buf19), .Y(random_clk_bf3__1661), );
  CLKBUF3 CLKBUF3__1662 (.Y(random_clk_bf3__1662), .A(clk_bF_buf19), );
  CLKBUF3 CLKBUF3__1681 (.A(clk_bF_buf10), .Y(random_clk_bf3__1681), );
  CLKBUF3 CLKBUF3__1682 (.Y(random_clk_bf3__1682), .A(clk_bF_buf10), );
  CLKBUF3 CLKBUF3__1701 (.A(clk_bF_buf1), .Y(random_clk_bf3__1701), );
  CLKBUF3 CLKBUF3__1702 (.Y(random_clk_bf3__1702), .A(clk_bF_buf1), );
  CLKBUF3 CLKBUF3__1721 (.A(clk_bF_buf90), .Y(random_clk_bf3__1721), );
  CLKBUF3 CLKBUF3__1722 (.Y(random_clk_bf3__1722), .A(clk_bF_buf90), );
  CLKBUF3 CLKBUF3__1741 (.A(clk_bF_buf81), .Y(random_clk_bf3__1741), );
  CLKBUF3 CLKBUF3__1742 (.Y(random_clk_bf3__1742), .A(clk_bF_buf81), );
  CLKBUF3 CLKBUF3__1761 (.A(clk_bF_buf72), .Y(random_clk_bf3__1761), );
  CLKBUF3 CLKBUF3__1762 (.Y(random_clk_bf3__1762), .A(clk_bF_buf72), );
  CLKBUF3 CLKBUF3__1781 (.A(clk_bF_buf63), .Y(random_clk_bf3__1781), );
  CLKBUF3 CLKBUF3__1782 (.Y(random_clk_bf3__1782), .A(clk_bF_buf63), );
  CLKBUF3 CLKBUF3__1801 (.A(clk_bF_buf54), .Y(random_clk_bf3__1801), );
  CLKBUF3 CLKBUF3__1802 (.Y(random_clk_bf3__1802), .A(clk_bF_buf54), );
  CLKBUF3 CLKBUF3__1821 (.A(clk_bF_buf45), .Y(random_clk_bf3__1821), );
  CLKBUF3 CLKBUF3__1822 (.Y(random_clk_bf3__1822), .A(clk_bF_buf45), );
  CLKBUF3 CLKBUF3__1841 (.A(clk_bF_buf36), .Y(random_clk_bf3__1841), );
  CLKBUF3 CLKBUF3__1842 (.Y(random_clk_bf3__1842), .A(clk_bF_buf36), );
  CLKBUF3 CLKBUF3__1861 (.A(clk_bF_buf27), .Y(random_clk_bf3__1861), );
  CLKBUF3 CLKBUF3__1862 (.Y(random_clk_bf3__1862), .A(clk_bF_buf27), );
  CLKBUF3 CLKBUF3__1881 (.A(clk_bF_buf18), .Y(random_clk_bf3__1881), );
  CLKBUF3 CLKBUF3__1882 (.Y(random_clk_bf3__1882), .A(clk_bF_buf18), );
  CLKBUF3 CLKBUF3__1901 (.A(clk_bF_buf9), .Y(random_clk_bf3__1901), );
  CLKBUF3 CLKBUF3__1902 (.Y(random_clk_bf3__1902), .A(clk_bF_buf9), );
  CLKBUF2 CLKBUF2__1 (.Y(clock_bf2__1), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__2 (.Y(clock_bf2__2), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__3 (.Y(clock_bf2__3), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__4 (.Y(clock_bf2__4), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__5 (.Y(clock_bf2__5), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__6 (.Y(clock_bf2__6), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__7 (.Y(clock_bf2__7), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__8 (.Y(clock_bf2__8), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__9 (.Y(clock_bf2__9), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__10 (.Y(clock_bf2__10), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__11 (.Y(clock_bf2__11), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__12 (.Y(clock_bf2__12), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__13 (.Y(clock_bf2__13), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__14 (.Y(clock_bf2__14), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__15 (.Y(clock_bf2__15), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__16 (.Y(clock_bf2__16), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__17 (.Y(clock_bf2__17), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__18 (.Y(clock_bf2__18), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__19 (.Y(clock_bf2__19), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__20 (.Y(clock_bf2__20), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__21 (.Y(clock_bf2__21), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__22 (.Y(clock_bf2__22), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__23 (.Y(clock_bf2__23), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__24 (.Y(clock_bf2__24), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__25 (.Y(clock_bf2__25), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__26 (.Y(clock_bf2__26), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__27 (.Y(clock_bf2__27), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__28 (.Y(clock_bf2__28), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__29 (.Y(clock_bf2__29), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__30 (.Y(clock_bf2__30), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__31 (.Y(clock_bf2__31), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__1 (.Y(clock_bf2__1), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__2 (.Y(clock_bf2__2), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__3 (.Y(clock_bf2__3), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__4 (.Y(clock_bf2__4), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__5 (.Y(clock_bf2__5), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__6 (.Y(clock_bf2__6), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__7 (.Y(clock_bf2__7), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__8 (.Y(clock_bf2__8), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__9 (.Y(clock_bf2__9), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__10 (.Y(clock_bf2__10), .A(clk_bF_buf98), );
  CLKBUF2 CLKBUF2__11 (.Y(clock_bf2__11), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__12 (.Y(clock_bf2__12), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__13 (.Y(clock_bf2__13), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__14 (.Y(clock_bf2__14), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__15 (.Y(clock_bf2__15), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__16 (.Y(clock_bf2__16), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__17 (.Y(clock_bf2__17), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__18 (.Y(clock_bf2__18), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__19 (.Y(clock_bf2__19), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__20 (.Y(clock_bf2__20), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__21 (.Y(clock_bf2__21), .A(clk_bF_buf97), );
  CLKBUF2 CLKBUF2__22 (.Y(clock_bf2__22), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__23 (.Y(clock_bf2__23), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__24 (.Y(clock_bf2__24), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__25 (.Y(clock_bf2__25), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__26 (.Y(clock_bf2__26), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__27 (.Y(clock_bf2__27), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__28 (.Y(clock_bf2__28), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__29 (.Y(clock_bf2__29), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__30 (.Y(clock_bf2__30), .A(clk_bF_buf0), );
  CLKBUF2 CLKBUF2__31 (.Y(clock_bf2__31), .A(clk_bF_buf0), );
endmodule

