module spi_slave ( gnd, vdd, SCK, SDI, CSB, idata, SDO, sdoenb, odata, oaddr, rdstb, wrstb);

input gnd, vdd;
input SCK;
input SDI;
input CSB;
output SDO;
output sdoenb;
output rdstb;
output wrstb;
input [7:0] idata;
output [7:0] odata;
output [7:0] oaddr;

CLKBUF1 CLKBUF1_1 ( .gnd(gnd), .vdd(vdd), .A(SCK), .Y(SCK_bF_buf4) );
CLKBUF1 CLKBUF1_2 ( .gnd(gnd), .vdd(vdd), .A(SCK), .Y(SCK_bF_buf3) );
CLKBUF1 CLKBUF1_3 ( .gnd(gnd), .vdd(vdd), .A(SCK), .Y(SCK_bF_buf2) );
CLKBUF1 CLKBUF1_4 ( .gnd(gnd), .vdd(vdd), .A(SCK), .Y(SCK_bF_buf1) );
CLKBUF1 CLKBUF1_5 ( .gnd(gnd), .vdd(vdd), .A(SCK), .Y(SCK_bF_buf0) );
BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_13__bF_buf5) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_13__bF_buf4) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_13__bF_buf3) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_13__bF_buf2) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_13__bF_buf1) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(_13__bF_buf0) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .Y(state_0_bF_buf3_) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .Y(state_0_bF_buf2_) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .Y(state_0_bF_buf1_) );
BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .Y(state_0_bF_buf0_) );
BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .Y(state_2_bF_buf3_) );
BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .Y(state_2_bF_buf2_) );
BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .Y(state_2_bF_buf1_) );
BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .Y(state_2_bF_buf0_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(addr_7_), .B(state_0_bF_buf3_), .Y(_157_) );
INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(state_0_bF_buf2_), .Y(_158_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(addr_6_), .Y(_159_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(state_2_bF_buf3_), .B(_159_), .Y(_160_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(addr_0_), .B(addr_1_), .Y(_161_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(addr_2_), .B(addr_3_), .Y(_15_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(addr_4_), .B(addr_5_), .Y(_16_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_15_), .C(_16_), .Y(_17_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(fixed_2_), .B(fixed_1_), .Y(_18_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(fixed_0_), .Y(_19_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(count_2_), .B(count_1_), .Y(_20_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(count_0_), .C(_20_), .Y(_21_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_19_), .C(_17_), .Y(_22_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(state_2_bF_buf2_), .B(_159_), .Y(_23_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(state_2_bF_buf1_), .B(addr_7_), .C(_23_), .Y(_24_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_160_), .B(_22_), .C(_24_), .Y(_25_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_160_), .Y(_26_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(addr_0_), .B(addr_1_), .Y(_27_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(addr_2_), .B(addr_3_), .Y(_28_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(addr_4_), .B(addr_5_), .Y(_29_) );
NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_28_), .C(_29_), .Y(_30_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(fixed_0_), .B(_18_), .Y(_31_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .Y(_32_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(count_2_), .B(count_0_), .C(count_1_), .Y(_33_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_33_), .Y(_34_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_34_), .C(_30_), .Y(_35_) );
NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(addr_7_), .B(_26_), .C(_35_), .Y(_36_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_36_), .C(_158_), .Y(_37_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_37_), .Y(_0__7_) );
INVX8 INVX8_2 ( .gnd(gnd), .vdd(vdd), .A(state_2_bF_buf0_), .Y(_38_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_32_), .Y(_39_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(state_0_bF_buf1_), .B(_38_), .Y(_40_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_164_), .C(_40_), .D(readmode), .Y(_41_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_39_), .C(_41_), .Y(_5_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(ldata_0_), .Y(_42_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(readmode), .B(state_1_), .Y(_7_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(count_0_), .Y(_43_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(count_1_), .Y(_44_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_44_), .Y(_45_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(count_2_), .B(_45_), .Y(_46_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(idata[0]), .B(_46_), .C(_7_), .Y(_47_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_7_), .C(_47_), .Y(_3__0_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(readmode), .Y(_48_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_32_), .C(ldata_1_), .Y(_49_) );
INVX8 INVX8_3 ( .gnd(gnd), .vdd(vdd), .A(_46_), .Y(_50_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_50_), .C(_7_), .Y(_51_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(idata[1]), .B(_50_), .C(_51_), .Y(_52_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_52_), .Y(_3__1_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(ldata_2_), .Y(_53_) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(idata[2]), .B(ldata_1_), .S(_46_), .Y(_54_) );
MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_54_), .S(_7_), .Y(_3__2_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_32_), .C(ldata_3_), .Y(_55_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_50_), .C(_7_), .Y(_56_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(idata[3]), .B(_50_), .C(_56_), .Y(_57_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(_57_), .Y(_3__3_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(ldata_4_), .Y(_58_) );
MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(idata[4]), .B(ldata_3_), .S(_46_), .Y(_59_) );
MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_59_), .S(_7_), .Y(_3__4_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_32_), .C(ldata_5_), .Y(_60_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_50_), .C(_7_), .Y(_61_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(idata[5]), .B(_50_), .C(_61_), .Y(_62_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_62_), .Y(_3__5_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(ldata_6_), .Y(_63_) );
MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(idata[6]), .B(ldata_5_), .S(_46_), .Y(_64_) );
MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_64_), .S(_7_), .Y(_3__6_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_32_), .C(ldata_7_), .Y(_65_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_50_), .C(_7_), .Y(_66_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(idata[7]), .B(_50_), .C(_66_), .Y(_67_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_67_), .Y(_3__7_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(_33_), .Y(_68_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(writemode), .C(_68_), .Y(_69_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_69_), .Y(_9_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(_68_), .C(_19_), .Y(_70_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_68_), .C(_70_), .Y(_10_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(state_2_bF_buf3_), .B(_33_), .Y(_71_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_33_), .C(_71_), .Y(_12_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_33_), .C(state_1_), .Y(_72_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_33_), .C(_72_), .Y(_11_) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(addr_0_), .Y(_73_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(state_2_bF_buf2_), .B(SDI), .Y(_74_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(state_2_bF_buf1_), .C(_74_), .Y(_162__0_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(addr_1_), .Y(_75_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(state_2_bF_buf0_), .B(addr_0_), .Y(_76_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(state_2_bF_buf3_), .C(_76_), .Y(_162__1_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(addr_2_), .B(_38_), .Y(_77_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_75_), .C(_77_), .Y(_162__2_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(addr_3_), .Y(_78_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(addr_2_), .Y(_79_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_79_), .Y(_80_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_80_), .Y(_81_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_78_), .B(state_2_bF_buf2_), .C(_81_), .Y(_162__3_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(addr_4_), .Y(_82_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(state_2_bF_buf1_), .B(addr_3_), .Y(_83_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(state_2_bF_buf0_), .C(_83_), .Y(_162__4_) );
INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(addr_5_), .Y(_84_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(state_2_bF_buf3_), .B(addr_4_), .Y(_85_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(state_2_bF_buf2_), .C(_85_), .Y(_162__5_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_84_), .C(_26_), .Y(_162__6_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_24_), .Y(_162__7_) );
INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(SDI), .Y(_86_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_163__1_), .Y(_87_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(state_2_bF_buf1_), .B(_32_), .Y(_88_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_88_), .Y(_89_) );
MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(_86_), .S(_89_), .Y(_4__0_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_163__2_), .Y(_90_) );
MUX2X1 MUX2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_87_), .S(_89_), .Y(_4__1_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_163__3_), .Y(_91_) );
MUX2X1 MUX2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_90_), .S(_89_), .Y(_4__2_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_163__4_), .Y(_92_) );
MUX2X1 MUX2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_92_), .B(_91_), .S(_89_), .Y(_4__3_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_163__5_), .Y(_93_) );
MUX2X1 MUX2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_92_), .S(_89_), .Y(_4__4_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_163__6_), .Y(_94_) );
MUX2X1 MUX2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_93_), .S(_89_), .Y(_4__5_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_163__7_), .Y(_95_) );
MUX2X1 MUX2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_94_), .S(_89_), .Y(_4__6_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(count_0_), .B(count_1_), .C(count_2_), .Y(_96_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(count_2_), .B(count_1_), .C(_96_), .Y(_97_) );
INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(_97_), .Y(_98_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_98_), .C(_158_), .Y(_99_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(fixed_0_), .B(_98_), .C(_99_), .Y(_100_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(fixed_2_), .B(fixed_1_), .C(_88_), .Y(_101_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_101_), .Y(_102_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(fixed_0_), .Y(_103_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(fixed_0_), .C(_158_), .Y(_104_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_104_), .C(_100_), .Y(_2__0_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(fixed_0_), .Y(_105_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_88_), .C(_68_), .Y(_106_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_106_), .B(fixed_1_), .Y(_107_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(fixed_2_), .B(_158_), .Y(_108_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(state_0_bF_buf0_), .B(_98_), .C(fixed_1_), .Y(_109_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(state_0_bF_buf3_), .B(_105_), .C(_98_), .Y(_110_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(state_0_bF_buf2_), .B(_106_), .C(_110_), .Y(_111_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_108_), .C(_111_), .D(_109_), .Y(_2__1_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(fixed_2_), .C(_107_), .Y(_112_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(fixed_2_), .B(_98_), .Y(_113_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(fixed_1_), .C(state_0_bF_buf1_), .Y(_114_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_114_), .C(_112_), .Y(_2__2_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(count_2_), .Y(_115_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(count_1_), .B(_43_), .Y(_116_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(state_0_bF_buf0_), .B(_115_), .C(_116_), .Y(_117_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(readmode), .B(_117_), .Y(_118_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_117_), .C(_118_), .Y(_6_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(state_0_bF_buf3_), .B(_46_), .Y(_119_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_158_), .C(writemode), .Y(_120_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_86_), .C(_120_), .Y(_8_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(state_0_bF_buf2_), .B(_39_), .Y(_121_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(count_0_), .Y(_1__0_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_43_), .C(_44_), .Y(_122_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_121_), .Y(_123_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(count_1_), .B(_123_), .Y(_124_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(_122_), .Y(_1__1_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_123_), .C(_124_), .D(_115_), .Y(_1__2_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_31_), .C(_34_), .Y(_125_) );
MUX2X1 MUX2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_162__0_), .B(_73_), .S(_125_), .Y(_126_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(state_0_bF_buf1_), .B(addr_0_), .Y(_127_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(state_0_bF_buf0_), .C(_127_), .Y(_0__0_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_21_), .Y(_128_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(state_0_bF_buf3_), .B(_73_), .Y(_129_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(state_2_bF_buf0_), .C(_129_), .Y(_130_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(state_0_bF_buf2_), .C(addr_1_), .Y(_131_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_131_), .Y(_0__1_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_34_), .Y(_132_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(addr_2_), .B(_161_), .Y(_133_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_133_), .Y(_134_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_27_), .C(_77_), .Y(_135_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_75_), .C(_158_), .Y(_136_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_135_), .C(_136_), .Y(_137_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(state_0_bF_buf1_), .B(_79_), .C(_137_), .Y(_0__2_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_132_), .Y(_138_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(state_2_bF_buf3_), .B(addr_3_), .Y(_139_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_138_), .C(_80_), .Y(_140_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_134_), .C(state_0_bF_buf0_), .Y(_141_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(state_0_bF_buf3_), .B(_140_), .C(_141_), .D(_78_), .Y(_0__3_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_28_), .Y(_142_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_31_), .C(_34_), .Y(_143_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(addr_4_), .Y(_144_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(addr_4_), .B(_143_), .Y(_145_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_145_), .C(_38_), .Y(_146_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(state_2_bF_buf2_), .B(addr_3_), .C(state_0_bF_buf2_), .Y(_147_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(state_0_bF_buf1_), .B(_82_), .C(_146_), .D(_147_), .Y(_0__4_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(addr_4_), .Y(_148_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_128_), .C(_84_), .Y(_149_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(addr_4_), .B(_142_), .Y(_150_) );
NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(addr_5_), .B(_150_), .C(_132_), .Y(_151_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_151_), .C(_38_), .Y(_152_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(state_2_bF_buf1_), .B(addr_4_), .C(state_0_bF_buf0_), .Y(_153_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(state_0_bF_buf3_), .B(_84_), .C(_152_), .D(_153_), .Y(_0__5_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(state_2_bF_buf0_), .B(addr_5_), .C(_35_), .D(_160_), .Y(_154_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(addr_6_), .B(state_2_bF_buf3_), .Y(_155_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_22_), .C(state_0_bF_buf2_), .Y(_156_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_159_), .B(state_0_bF_buf1_), .C(_156_), .D(_154_), .Y(_0__6_) );
INVX4 INVX4_3 ( .gnd(gnd), .vdd(vdd), .A(SCK_bF_buf4), .Y(_14_) );
INVX8 INVX8_4 ( .gnd(gnd), .vdd(vdd), .A(CSB), .Y(_13_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(ldata_7_), .Y(SDO) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_162__0_), .Y(oaddr[0]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_162__1_), .Y(oaddr[1]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_162__2_), .Y(oaddr[2]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_162__3_), .Y(oaddr[3]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_162__4_), .Y(oaddr[4]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_162__5_), .Y(oaddr[5]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_162__6_), .Y(oaddr[6]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_162__7_), .Y(oaddr[7]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(SDI), .Y(odata[0]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_163__1_), .Y(odata[1]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_163__2_), .Y(odata[2]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_163__3_), .Y(odata[3]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_163__4_), .Y(odata[4]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_163__5_), .Y(odata[5]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_163__6_), .Y(odata[6]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_163__7_), .Y(odata[7]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_164_), .Y(rdstb) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_165_), .Y(sdoenb) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_166_), .Y(wrstb) );
DFFSR DFFSR_1 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf3), .D(_5_), .Q(_164_), .R(_13__bF_buf5), .S(vdd) );
DFFSR DFFSR_2 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf2), .D(_10_), .Q(state_0_), .R(vdd), .S(_13__bF_buf4) );
DFFSR DFFSR_3 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf1), .D(_11_), .Q(state_1_), .R(_13__bF_buf3), .S(vdd) );
DFFSR DFFSR_4 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf0), .D(_12_), .Q(state_2_), .R(_13__bF_buf2), .S(vdd) );
DFFSR DFFSR_5 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf4), .D(_0__0_), .Q(addr_0_), .R(_13__bF_buf1), .S(vdd) );
DFFSR DFFSR_6 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf3), .D(_0__1_), .Q(addr_1_), .R(_13__bF_buf0), .S(vdd) );
DFFSR DFFSR_7 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf2), .D(_0__2_), .Q(addr_2_), .R(_13__bF_buf5), .S(vdd) );
DFFSR DFFSR_8 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf1), .D(_0__3_), .Q(addr_3_), .R(_13__bF_buf4), .S(vdd) );
DFFSR DFFSR_9 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf0), .D(_0__4_), .Q(addr_4_), .R(_13__bF_buf3), .S(vdd) );
DFFSR DFFSR_10 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf4), .D(_0__5_), .Q(addr_5_), .R(_13__bF_buf2), .S(vdd) );
DFFSR DFFSR_11 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf3), .D(_0__6_), .Q(addr_6_), .R(_13__bF_buf1), .S(vdd) );
DFFSR DFFSR_12 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf2), .D(_0__7_), .Q(addr_7_), .R(_13__bF_buf0), .S(vdd) );
DFFSR DFFSR_13 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf1), .D(_1__0_), .Q(count_0_), .R(_13__bF_buf5), .S(vdd) );
DFFSR DFFSR_14 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf0), .D(_1__1_), .Q(count_1_), .R(_13__bF_buf4), .S(vdd) );
DFFSR DFFSR_15 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf4), .D(_1__2_), .Q(count_2_), .R(_13__bF_buf3), .S(vdd) );
DFFSR DFFSR_16 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf3), .D(_8_), .Q(writemode), .R(_13__bF_buf2), .S(vdd) );
DFFSR DFFSR_17 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf2), .D(_6_), .Q(readmode), .R(_13__bF_buf1), .S(vdd) );
DFFSR DFFSR_18 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf1), .D(_2__0_), .Q(fixed_0_), .R(_13__bF_buf0), .S(vdd) );
DFFSR DFFSR_19 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf0), .D(_2__1_), .Q(fixed_1_), .R(_13__bF_buf5), .S(vdd) );
DFFSR DFFSR_20 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf4), .D(_2__2_), .Q(fixed_2_), .R(_13__bF_buf4), .S(vdd) );
DFFSR DFFSR_21 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf3), .D(_4__0_), .Q(_163__1_), .R(_13__bF_buf3), .S(vdd) );
DFFSR DFFSR_22 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf2), .D(_4__1_), .Q(_163__2_), .R(_13__bF_buf2), .S(vdd) );
DFFSR DFFSR_23 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf1), .D(_4__2_), .Q(_163__3_), .R(_13__bF_buf1), .S(vdd) );
DFFSR DFFSR_24 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf0), .D(_4__3_), .Q(_163__4_), .R(_13__bF_buf0), .S(vdd) );
DFFSR DFFSR_25 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf4), .D(_4__4_), .Q(_163__5_), .R(_13__bF_buf5), .S(vdd) );
DFFSR DFFSR_26 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf3), .D(_4__5_), .Q(_163__6_), .R(_13__bF_buf4), .S(vdd) );
DFFSR DFFSR_27 ( .gnd(gnd), .vdd(vdd), .CLK(SCK_bF_buf2), .D(_4__6_), .Q(_163__7_), .R(_13__bF_buf3), .S(vdd) );
DFFSR DFFSR_28 ( .gnd(gnd), .vdd(vdd), .CLK(_14_), .D(_7_), .Q(_165_), .R(vdd), .S(_13__bF_buf2) );
DFFSR DFFSR_29 ( .gnd(gnd), .vdd(vdd), .CLK(_14_), .D(_9_), .Q(_166_), .R(_13__bF_buf1), .S(vdd) );
DFFSR DFFSR_30 ( .gnd(gnd), .vdd(vdd), .CLK(_14_), .D(_3__0_), .Q(ldata_0_), .R(_13__bF_buf0), .S(vdd) );
DFFSR DFFSR_31 ( .gnd(gnd), .vdd(vdd), .CLK(_14_), .D(_3__1_), .Q(ldata_1_), .R(_13__bF_buf5), .S(vdd) );
DFFSR DFFSR_32 ( .gnd(gnd), .vdd(vdd), .CLK(_14_), .D(_3__2_), .Q(ldata_2_), .R(_13__bF_buf4), .S(vdd) );
DFFSR DFFSR_33 ( .gnd(gnd), .vdd(vdd), .CLK(_14_), .D(_3__3_), .Q(ldata_3_), .R(_13__bF_buf3), .S(vdd) );
DFFSR DFFSR_34 ( .gnd(gnd), .vdd(vdd), .CLK(_14_), .D(_3__4_), .Q(ldata_4_), .R(_13__bF_buf2), .S(vdd) );
DFFSR DFFSR_35 ( .gnd(gnd), .vdd(vdd), .CLK(_14_), .D(_3__5_), .Q(ldata_5_), .R(_13__bF_buf1), .S(vdd) );
DFFSR DFFSR_36 ( .gnd(gnd), .vdd(vdd), .CLK(_14_), .D(_3__6_), .Q(ldata_6_), .R(_13__bF_buf0), .S(vdd) );
DFFSR DFFSR_37 ( .gnd(gnd), .vdd(vdd), .CLK(_14_), .D(_3__7_), .Q(ldata_7_), .R(_13__bF_buf5), .S(vdd) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(SDI), .Y(_163__0_) );
endmodule
