module add ( gnd, vdd, a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, rst, on, clk, out);

input gnd, vdd;
input a;
input b;
input c;
input d;
input e;
input f;
input g;
input h;
input i;
input j;
input k;
input l;
input m;
input n;
input o;
input p;
input q;
input r;
input s;
input t;
input u;
input v;
input w;
input x;
input y;
input rst;
input on;
input clk;
output out;

NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(g), .B(_24_), .Y(_25_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(g), .Y(_26_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_23_), .C(_26_), .D(_25_), .Y(_27_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_23_), .Y(_28_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(g), .Y(_29_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_28_), .Y(_30_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_27_), .C(_30_), .Y(_31_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_11_), .Y(_32_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_28_), .Y(_33_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(g), .Y(_34_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_23_), .C(_34_), .Y(_35_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_35_), .C(_32_), .Y(_36_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(j), .B(b), .Y(_37_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_37_), .Y(_38_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_36_), .C(_38_), .Y(_39_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_32_), .C(_35_), .Y(_40_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_27_), .C(_16_), .Y(_41_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_40_), .C(_41_), .Y(_42_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(a), .B(h), .Y(_43_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(a), .B(h), .Y(_44_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(_44_), .Y(_45_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_43_), .Y(_46_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(q), .Y(_47_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(f), .B(y), .Y(_48_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_48_), .Y(_49_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(f), .Y(_50_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(y), .B(_50_), .Y(_51_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(y), .Y(_52_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(f), .B(_52_), .Y(_53_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_51_), .B(_53_), .C(q), .Y(_54_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_54_), .C(_46_), .Y(_55_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_45_), .Y(_56_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(q), .B(_51_), .C(_53_), .Y(_57_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_48_), .Y(_58_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_57_), .C(_58_), .Y(_59_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(c), .B(k), .Y(_60_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(l), .Y(_61_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_61_), .Y(_62_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(_59_), .C(_62_), .Y(_63_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_58_), .C(_56_), .Y(_64_) );
NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_54_), .C(_49_), .Y(_65_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_64_), .C(_61_), .Y(_66_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(d), .B(_66_), .C(_63_), .Y(_67_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(d), .Y(_68_) );
NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_61_), .C(_65_), .Y(_69_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(_55_), .C(_62_), .Y(_70_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_70_), .C(_68_), .Y(_71_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_67_), .B(_71_), .C(_39_), .D(_42_), .Y(_72_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_41_), .C(_37_), .Y(_73_) );
NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_38_), .C(_31_), .Y(_74_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_67_), .B(_71_), .Y(_75_) );
NOR3X1 NOR3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_74_), .C(_75_), .Y(_1_) );
NOR3X1 NOR3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_2_), .B(_72_), .C(_1_), .Y(_0_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_76_), .Y(out) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(_0_), .Q(_76_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(_2_) );
XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(v), .B(t), .Y(_3_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(x), .B(n), .Y(_4_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(x), .B(n), .Y(_5_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_5_), .C(s), .Y(_6_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(s), .Y(_7_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(x), .B(n), .Y(_8_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(x), .B(n), .Y(_9_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_8_), .C(_9_), .Y(_10_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_3_), .B(_6_), .C(_10_), .Y(_11_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_3_), .Y(_12_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_9_), .C(_7_), .Y(_13_) );
NOR3X1 NOR3X1_7 ( .gnd(gnd), .vdd(vdd), .A(s), .B(_5_), .C(_4_), .Y(_14_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_13_), .C(_12_), .Y(_15_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_15_), .Y(_16_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(o), .B(m), .Y(_17_) );
XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(e), .B(r), .Y(_18_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_17_), .Y(_19_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(o), .B(m), .Y(_20_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(o), .B(m), .Y(_21_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(e), .B(r), .Y(_22_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .C(_22_), .Y(_23_) );
XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(w), .B(u), .Y(_24_) );
endmodule
