`ifndef _TIMESCALE_VH_
	`timescale 1ns/1ps
`endif
