module map9v3 ( gnd, vdd, clock, reset, start, N, dp, done, counter, sr);

input gnd;
input vdd;
input clock;
input reset;
input start;
output done;
input [3:0] N;
output [3:0] dp;
output [2:0] counter;
output [2:0] sr;

CLKBUF1 CLKBUF1_1 ( .gnd(gnd), .vdd(vdd), .A(clock), .Y(clock_bF_buf3) );
CLKBUF1 CLKBUF1_2 ( .gnd(gnd), .vdd(vdd), .A(clock), .Y(clock_bF_buf2) );
CLKBUF1 CLKBUF1_3 ( .gnd(gnd), .vdd(vdd), .A(clock), .Y(clock_bF_buf1) );
CLKBUF1 CLKBUF1_4 ( .gnd(gnd), .vdd(vdd), .A(clock), .Y(clock_bF_buf0) );
BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(_8_), .Y(_8__bF_buf3) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(_8_), .Y(_8__bF_buf2) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(_8_), .Y(_8__bF_buf1) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(_8_), .Y(_8__bF_buf0) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_44__1_), .Y(counter[1]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_44__2_), .Y(counter[2]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_45_), .Y(done) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_46__0_), .Y(dp[0]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_46__1_), .Y(dp[1]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_46__2_), .Y(dp[2]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_46__3_), .Y(dp[3]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_47__0_), .Y(sr[0]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_47__1_), .Y(sr[1]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_47__2_), .Y(sr[2]) );
DFFSR DFFSR_1 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf0), .D(_4_), .Q(state_0_), .R(vdd), .S(_8__bF_buf2) );
DFFSR DFFSR_2 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf2), .D(_6_), .Q(state_1_), .R(_8__bF_buf0), .S(vdd) );
DFFSR DFFSR_3 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf2), .D(_5_), .Q(state_2_), .R(_8__bF_buf1), .S(vdd) );
DFFSR DFFSR_4 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf1), .D(_7_), .Q(state_3_), .R(_8__bF_buf1), .S(vdd) );
DFFSR DFFSR_5 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf1), .D(state_2_), .Q(state_4_), .R(_8__bF_buf0), .S(vdd) );
DFFSR DFFSR_6 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf2), .D(start), .Q(startbuf_0_), .R(_8__bF_buf0), .S(vdd) );
DFFSR DFFSR_7 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf2), .D(startbuf_0_), .Q(startbuf_1_), .R(_8__bF_buf2), .S(vdd) );
DFFSR DFFSR_8 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf3), .D(_0__0_), .Q(_44__0_), .R(_8__bF_buf3), .S(vdd) );
DFFSR DFFSR_9 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf1), .D(_0__1_), .Q(_44__1_), .R(_8__bF_buf1), .S(vdd) );
DFFSR DFFSR_10 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf1), .D(_0__2_), .Q(_44__2_), .R(_8__bF_buf1), .S(vdd) );
DFFSR DFFSR_11 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf3), .D(_3__0_), .Q(_47__0_), .R(_8__bF_buf3), .S(vdd) );
DFFSR DFFSR_12 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf3), .D(_3__1_), .Q(_47__1_), .R(_8__bF_buf3), .S(vdd) );
DFFSR DFFSR_13 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf3), .D(_3__2_), .Q(_47__2_), .R(_8__bF_buf3), .S(vdd) );
DFFSR DFFSR_14 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf0), .D(_2__0_), .Q(_46__0_), .R(_8__bF_buf2), .S(vdd) );
DFFSR DFFSR_15 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf3), .D(_2__1_), .Q(_46__1_), .R(_8__bF_buf3), .S(vdd) );
DFFSR DFFSR_16 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf0), .D(_2__2_), .Q(_46__2_), .R(_8__bF_buf2), .S(vdd) );
DFFSR DFFSR_17 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf0), .D(_2__3_), .Q(_46__3_), .R(_8__bF_buf2), .S(vdd) );
DFFSR DFFSR_18 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf2), .D(_1_), .Q(_45_), .R(_8__bF_buf0), .S(vdd) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .Y(_9_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .Y(_10_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_44__1_), .B(_44__0_), .C(_44__2_), .Y(_11_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_10_), .C(_9_), .Y(_7_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .Y(_12_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .Y(_13_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(startbuf_0_), .Y(_14_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(startbuf_1_), .B(_14_), .Y(_15_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_12_), .C(_13_), .Y(_6_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_46__1_), .Y(_16_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_47__0_), .Y(_17_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(_9_), .C(_10_), .Y(_18_) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_17_), .S(_18_), .Y(_2__1_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_46__2_), .Y(_19_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_47__1_), .Y(_20_) );
MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_20_), .S(_18_), .Y(_2__2_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_46__3_), .Y(_21_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_47__2_), .Y(_22_) );
MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_22_), .S(_18_), .Y(_2__3_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_46__0_), .Y(_23_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(N[0]), .Y(_24_) );
MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_24_), .S(_18_), .Y(_2__0_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .B(_47__1_), .Y(_25_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .B(_47__0_), .C(_25_), .Y(_26_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(_26_), .Y(_3__0_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(state_3_), .C(_25_), .Y(_27_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_9_), .Y(_3__2_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_47__0_), .C(_9_), .Y(_28_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_20_), .C(_28_), .Y(_3__1_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_45_), .Y(_29_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .Y(_30_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .B(_10_), .C(_30_), .Y(_31_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_31_), .C(state_0_), .Y(_1_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_44__0_), .B(_10_), .Y(_32_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_44__0_), .Y(_33_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .B(_33_), .C(state_0_), .Y(_34_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(N[1]), .C(_34_), .D(_32_), .Y(_0__0_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .B(_44__1_), .C(_33_), .Y(_35_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_44__1_), .Y(_36_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_44__0_), .C(_36_), .Y(_37_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_35_), .C(_37_), .Y(_38_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(N[2]), .Y(_39_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_38_), .Y(_0__1_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(N[2]), .B(N[3]), .Y(_40_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_44__1_), .B(_44__0_), .Y(_41_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(_10_), .C(_44__2_), .Y(_42_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .B(_11_), .C(state_0_), .Y(_43_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(_40_), .C(_43_), .D(_42_), .Y(_0__2_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(state_1_), .Y(_4_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(state_3_), .Y(_5_) );
INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(_8_) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_44__0_), .Y(counter[0]) );
endmodule
