module divider ( gnd, vdd, clk, sign, start, dividend, divider, quotient, remainder, ready);

input gnd, vdd;
input clk;
input sign;
input start;
output ready;
input [3:0] dividend;
input [3:0] divider;
output [3:0] quotient;
output [3:0] remainder;

CLKBUF1 CLKBUF1_1 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf4) );
CLKBUF1 CLKBUF1_2 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf3) );
CLKBUF1 CLKBUF1_3 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf2) );
CLKBUF1 CLKBUF1_4 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf1) );
CLKBUF1 CLKBUF1_5 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf0) );
BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(_65_), .Y(_65__bF_buf3) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(_65_), .Y(_65__bF_buf2) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(_65_), .Y(_65__bF_buf1) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(_65_), .Y(_65__bF_buf0) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(_181_), .Y(_181__bF_buf3) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(_181_), .Y(_181__bF_buf2) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(_181_), .Y(_181__bF_buf1) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(_181_), .Y(_181__bF_buf0) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_22_), .Y(_23_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_4_), .Y(_24_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(dividend_copy_4_), .Y(_25_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_4_), .B(_24_), .Y(_26_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_25_), .Y(_27_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_23_), .Y(_28_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_5_), .B(_21_), .C(_25_), .Y(_29_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(divider_copy_5_), .C(_29_), .Y(_30_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_18_), .C(_30_), .Y(_31_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_6_), .B(_182_), .Y(_32_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_32_), .C(_7_), .Y(_33_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_7_), .B(dividend_copy_7_), .Y(_34_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_33_), .Y(_35_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_1_), .Y(_36_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_1_), .B(_36_), .Y(_37_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_0_), .B(_180_), .Y(_38_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_1_), .B(_36_), .Y(_39_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_39_), .C(_37_), .Y(_40_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_3_), .B(divider_copy_3_), .Y(_41_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_2_), .B(divider_copy_2_), .Y(_42_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(_42_), .Y(_43_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_3_), .Y(_44_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_3_), .B(_44_), .Y(_45_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_2_), .Y(_46_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_2_), .B(_46_), .Y(_47_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(_47_), .C(_45_), .Y(_48_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_43_), .C(_48_), .Y(_49_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_27_), .Y(_50_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(_51_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_50_), .C(_51_), .Y(_52_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_6_), .B(divider_copy_6_), .Y(_53_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_52_), .Y(_54_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_34_), .Y(_55_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_54_), .C(_55_), .Y(_56_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_56_), .C(_181__bF_buf0), .Y(_57_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_180_), .C(dividend_copy_0_), .Y(_58_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(_57_), .Y(_59_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_59_), .C(start), .Y(_60_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(start), .C(_60_), .D(_58_), .Y(_2__0_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(dividend[1]), .Y(_61_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(dividend[3]), .B(sign), .Y(_62_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_62_), .Y(_63_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(dividend[0]), .B(_63_), .Y(_64_) );
INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(start), .Y(_65_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_64_), .C(_65__bF_buf2), .Y(_66_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_64_), .C(_66_), .Y(_67_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_9_), .C(_10_), .Y(_68_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_39_), .C(_38_), .Y(_69_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_69_), .C(_57_), .Y(_70_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(dividend_copy_1_), .C(_65__bF_buf3), .Y(_71_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_70_), .C(_67_), .Y(_2__1_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_61_), .C(_62_), .Y(_72_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(dividend[2]), .B(_72_), .C(_65__bF_buf2), .Y(_73_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(dividend[2]), .B(_72_), .C(_73_), .Y(_74_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_35_), .Y(_75_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_1_), .C(_177_), .Y(_76_) );
XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_13_), .Y(_77_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_77_), .C(_76_), .Y(_78_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_78_), .B(start), .C(_74_), .Y(_2__2_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_61_), .Y(_79_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(dividend[2]), .C(sign), .Y(_80_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(dividend[3]), .B(start), .C(_80_), .Y(_81_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_42_), .C(_47_), .Y(_82_) );
XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_41_), .Y(_83_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_57_), .Y(_84_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(dividend_copy_3_), .C(_65__bF_buf3), .Y(_85_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_84_), .C(_81_), .Y(_2__3_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_27_), .Y(_86_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_18_), .Y(_87_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(_86_), .Y(_88_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_59_), .Y(_89_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_1_), .C(dividend_copy_4_), .Y(_90_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_89_), .C(start), .Y(_2__4_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_86_), .Y(_91_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_23_), .Y(_92_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(dividend_copy_5_), .C(_65__bF_buf0), .Y(_93_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(_92_), .C(_93_), .Y(_2__5_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_53_), .Y(_94_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_94_), .C(_59_), .Y(_95_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_1_), .C(dividend_copy_6_), .Y(_96_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(_95_), .C(start), .Y(_2__6_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_1_), .C(dividend_copy_7_), .Y(_97_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(start), .B(_97_), .Y(_2__7_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(dividend[3]), .B(divider[3]), .Y(_98_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(sign), .B(divider[3]), .Y(_99_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_99_), .Y(_100_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_100_), .C(_98_), .Y(_101_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(negative_output), .B(_65__bF_buf2), .Y(_102_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_65__bF_buf2), .C(_102_), .Y(_4_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_181__bF_buf0), .B(divider_copy_0_), .C(_65__bF_buf3), .Y(_103_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_181__bF_buf0), .C(_103_), .Y(_3__0_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_181__bF_buf2), .B(divider_copy_1_), .C(_65__bF_buf3), .Y(_104_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_181__bF_buf2), .C(_104_), .Y(_3__1_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_181__bF_buf2), .B(divider_copy_2_), .C(_65__bF_buf3), .Y(_105_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_181__bF_buf2), .C(_105_), .Y(_3__2_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(bit_5_), .C(_24_), .Y(_106_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_181__bF_buf2), .B(divider_copy_3_), .C(_106_), .Y(_107_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(start), .B(divider[0]), .Y(_108_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(start), .C(_108_), .Y(_3__3_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_5_), .B(_1_), .Y(_109_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_181__bF_buf1), .B(divider_copy_4_), .C(_65__bF_buf0), .Y(_110_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(divider[1]), .Y(_111_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(divider[0]), .B(_100_), .Y(_112_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_112_), .C(_65__bF_buf0), .Y(_113_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_112_), .C(_113_), .Y(_114_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_109_), .C(_114_), .Y(_3__4_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_6_), .B(_1_), .Y(_115_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_181__bF_buf1), .B(divider_copy_5_), .C(_65__bF_buf0), .Y(_116_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(divider[0]), .Y(_117_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_111_), .C(_99_), .Y(_118_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(divider[2]), .B(_118_), .C(_65__bF_buf2), .Y(_119_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(divider[2]), .B(_118_), .C(_119_), .Y(_120_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(_115_), .C(_120_), .Y(_3__5_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_1_), .Y(_121_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_7_), .B(_1_), .C(_121_), .Y(_122_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_111_), .Y(_123_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_123_), .B(divider[2]), .C(sign), .Y(_124_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(divider[3]), .B(_124_), .C(_65__bF_buf2), .Y(_125_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_65__bF_buf0), .B(_122_), .C(_125_), .Y(_3__6_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_7_), .B(_65__bF_buf0), .Y(_126_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_181__bF_buf1), .Y(_3__7_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(bit_5_), .C(_65__bF_buf1), .Y(_127_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(bit_0_), .Y(_128_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_128_), .Y(_0__0_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_127_), .Y(_129_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(bit_1_), .B(bit_0_), .Y(_130_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_130_), .C(_129_), .Y(_131_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_131_), .Y(_0__1_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(bit_1_), .B(bit_0_), .C(bit_2_), .Y(_132_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_132_), .Y(_133_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1_), .B(_133_), .C(_65__bF_buf1), .Y(_0__2_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(bit_2_), .C(bit_3_), .Y(_134_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(_134_), .C(_127_), .Y(_0__3_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(bit_5_), .B(_65__bF_buf1), .Y(_135_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(bit_3_), .C(bit_4_), .Y(_136_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(start), .B(_136_), .C(_169_), .D(_135_), .Y(_0__4_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(bit_4_), .C(bit_5_), .Y(_137_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(start), .B(_137_), .Y(_0__5_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(quotient_temp_0_), .Y(_138_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_181__bF_buf0), .C(_57_), .Y(_139_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_65__bF_buf3), .Y(_6__0_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(bit_5_), .C(_138_), .Y(_140_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_181__bF_buf3), .B(quotient_temp_1_), .C(_140_), .Y(_141_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(start), .B(_141_), .Y(_6__1_) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(quotient_temp_1_), .Y(_142_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_181__bF_buf3), .B(quotient_temp_2_), .C(_65__bF_buf1), .Y(_143_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_181__bF_buf3), .C(_143_), .Y(_6__2_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_183__0_), .B(_1_), .Y(_144_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_57_), .C(start), .Y(_5__0_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_138_), .Y(_145_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_56_), .C(negative_output), .Y(_146_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_146_), .Y(_147_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_183__1_), .Y(_148_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(start), .B(_148_), .C(_127_), .Y(_149_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_140_), .C(_149_), .Y(_150_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(_145_), .C(_150_), .Y(_5__1_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_55_), .C(_54_), .Y(_151_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_33_), .Y(_152_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_152_), .C(_151_), .Y(_153_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(negative_output), .B(_153_), .Y(_154_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(quotient_temp_1_), .B(_1_), .C(_154_), .Y(_155_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_138_), .C(_146_), .Y(_156_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_1_), .C(_156_), .Y(_157_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_181__bF_buf3), .B(_183__2_), .C(_65__bF_buf1), .Y(_158_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_157_), .C(_158_), .Y(_5__2_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(quotient_temp_2_), .Y(_159_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_142_), .Y(_160_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_160_), .C(_159_), .Y(_161_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(quotient_temp_1_), .C(negative_output), .Y(_162_) );
AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(quotient_temp_2_), .B(_162_), .C(_1_), .Y(_163_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_181__bF_buf3), .B(_183__3_), .C(_65__bF_buf1), .Y(_164_) );
AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_163_), .C(_164_), .Y(_5__3_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(del_ready), .B(_181__bF_buf1), .Y(_184_) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_0_), .Y(remainder[0]) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(bit_1_), .B(bit_0_), .Y(_165_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_165_), .Y(_166_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(bit_2_), .Y(_167_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(bit_3_), .Y(_168_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(bit_4_), .Y(_169_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(bit_5_), .B(_169_), .Y(_1_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_1_), .Y(_170_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_0_), .Y(_171_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_0_), .B(dividend_copy_1_), .C(negative_output), .Y(_172_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_172_), .Y(_173_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_170_), .C(_173_), .Y(_174_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(negative_output), .B(_170_), .C(_174_), .Y(_185__1_) );
XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(dividend_copy_2_), .Y(_185__2_) );
INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_3_), .Y(_175_) );
INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(negative_output), .Y(_176_) );
INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_2_), .Y(_177_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_177_), .C(_172_), .Y(_178_) );
XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_175_), .Y(_185__3_) );
INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(dividend[0]), .Y(_179_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_0_), .Y(_180_) );
INVX8 INVX8_2 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(_181_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_6_), .Y(_182_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_6_), .B(_182_), .Y(_7_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_1_), .B(_170_), .Y(_8_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_0_), .B(_171_), .Y(_9_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_1_), .B(_170_), .Y(_10_) );
AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_10_), .C(_8_), .Y(_11_) );
XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_3_), .B(divider_copy_3_), .Y(_12_) );
XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_2_), .B(divider_copy_2_), .Y(_13_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_13_), .Y(_14_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_3_), .B(_175_), .Y(_15_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_2_), .B(_177_), .Y(_16_) );
AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_12_), .C(_15_), .Y(_17_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_11_), .C(_17_), .Y(_18_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_5_), .Y(_19_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_5_), .B(_19_), .Y(_20_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(divider_copy_5_), .Y(_21_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(dividend_copy_5_), .B(_21_), .Y(_22_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_183__0_), .Y(quotient[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_183__1_), .Y(quotient[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_183__2_), .Y(quotient[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_183__3_), .Y(quotient[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_184_), .Y(ready) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_185__1_), .Y(remainder[1]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_185__2_), .Y(remainder[2]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_185__3_), .Y(remainder[3]) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_6__0_), .Q(quotient_temp_0_) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_6__1_), .Q(quotient_temp_1_) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_6__2_), .Q(quotient_temp_2_) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_2__0_), .Q(dividend_copy_0_) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_2__1_), .Q(dividend_copy_1_) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_2__2_), .Q(dividend_copy_2_) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_2__3_), .Q(dividend_copy_3_) );
DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_2__4_), .Q(dividend_copy_4_) );
DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_2__5_), .Q(dividend_copy_5_) );
DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_2__6_), .Q(dividend_copy_6_) );
DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_2__7_), .Q(dividend_copy_7_) );
DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_5__0_), .Q(_183__0_) );
DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_5__1_), .Q(_183__1_) );
DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_5__2_), .Q(_183__2_) );
DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_5__3_), .Q(_183__3_) );
DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_3__0_), .Q(divider_copy_0_) );
DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_3__1_), .Q(divider_copy_1_) );
DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_3__2_), .Q(divider_copy_2_) );
DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_3__3_), .Q(divider_copy_3_) );
DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_3__4_), .Q(divider_copy_4_) );
DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_3__5_), .Q(divider_copy_5_) );
DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3__6_), .Q(divider_copy_6_) );
DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3__7_), .Q(divider_copy_7_) );
DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_4_), .Q(negative_output) );
DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0__0_), .Q(bit_0_) );
DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0__1_), .Q(bit_1_) );
DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0__2_), .Q(bit_2_) );
DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0__3_), .Q(bit_3_) );
DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0__4_), .Q(bit_4_) );
DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__5_), .Q(bit_5_) );
DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_1_), .Q(del_ready) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(remainder[0]), .Y(_185__0_) );
endmodule
