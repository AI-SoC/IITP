module picorv32_regs ( gnd, vdd, clk, wen, waddr, raddr1, raddr2, wdata, rdata1, rdata2);

input gnd, vdd;
input clk;
input wen;
input [5:0] waddr;
input [5:0] raddr1;
input [5:0] raddr2;
input [31:0] wdata;
output [31:0] rdata1;
output [31:0] rdata2;

BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(raddr2_1_bF_buf14_), .Y(raddr2_1_bF_buf14_bF_buf3_) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(raddr2_1_bF_buf14_), .Y(raddr2_1_bF_buf14_bF_buf2_) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(raddr2_1_bF_buf14_), .Y(raddr2_1_bF_buf14_bF_buf1_) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(raddr2_1_bF_buf14_), .Y(raddr2_1_bF_buf14_bF_buf0_) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf8) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf7) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf6) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf5) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf4) );
BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf3) );
BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf2) );
BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf1) );
BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf0) );
BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf13_), .Y(raddr1_1_bF_buf13_bF_buf3_) );
BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf13_), .Y(raddr1_1_bF_buf13_bF_buf2_) );
BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf13_), .Y(raddr1_1_bF_buf13_bF_buf1_) );
BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf13_), .Y(raddr1_1_bF_buf13_bF_buf0_) );
BUFX4 BUFX4_18 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf10_), .Y(raddr1_1_bF_buf10_bF_buf3_) );
BUFX4 BUFX4_19 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf10_), .Y(raddr1_1_bF_buf10_bF_buf2_) );
BUFX4 BUFX4_20 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf10_), .Y(raddr1_1_bF_buf10_bF_buf1_) );
BUFX4 BUFX4_21 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf10_), .Y(raddr1_1_bF_buf10_bF_buf0_) );
BUFX4 BUFX4_22 ( .gnd(gnd), .vdd(vdd), .A(raddr2[0]), .Y(raddr2_0__hier0_bF_buf8) );
BUFX4 BUFX4_23 ( .gnd(gnd), .vdd(vdd), .A(raddr2[0]), .Y(raddr2_0__hier0_bF_buf7) );
BUFX4 BUFX4_24 ( .gnd(gnd), .vdd(vdd), .A(raddr2[0]), .Y(raddr2_0__hier0_bF_buf6) );
BUFX4 BUFX4_25 ( .gnd(gnd), .vdd(vdd), .A(raddr2[0]), .Y(raddr2_0__hier0_bF_buf5) );
BUFX4 BUFX4_26 ( .gnd(gnd), .vdd(vdd), .A(raddr2[0]), .Y(raddr2_0__hier0_bF_buf4) );
BUFX4 BUFX4_27 ( .gnd(gnd), .vdd(vdd), .A(raddr2[0]), .Y(raddr2_0__hier0_bF_buf3) );
BUFX4 BUFX4_28 ( .gnd(gnd), .vdd(vdd), .A(raddr2[0]), .Y(raddr2_0__hier0_bF_buf2) );
BUFX4 BUFX4_29 ( .gnd(gnd), .vdd(vdd), .A(raddr2[0]), .Y(raddr2_0__hier0_bF_buf1) );
BUFX4 BUFX4_30 ( .gnd(gnd), .vdd(vdd), .A(raddr2[0]), .Y(raddr2_0__hier0_bF_buf0) );
BUFX4 BUFX4_31 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf9_), .Y(raddr1_1_bF_buf9_bF_buf3_) );
BUFX4 BUFX4_32 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf9_), .Y(raddr1_1_bF_buf9_bF_buf2_) );
BUFX4 BUFX4_33 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf9_), .Y(raddr1_1_bF_buf9_bF_buf1_) );
BUFX4 BUFX4_34 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf9_), .Y(raddr1_1_bF_buf9_bF_buf0_) );
BUFX4 BUFX4_35 ( .gnd(gnd), .vdd(vdd), .A(raddr1[0]), .Y(raddr1_0__hier0_bF_buf8) );
BUFX4 BUFX4_36 ( .gnd(gnd), .vdd(vdd), .A(raddr1[0]), .Y(raddr1_0__hier0_bF_buf7) );
BUFX4 BUFX4_37 ( .gnd(gnd), .vdd(vdd), .A(raddr1[0]), .Y(raddr1_0__hier0_bF_buf6) );
BUFX4 BUFX4_38 ( .gnd(gnd), .vdd(vdd), .A(raddr1[0]), .Y(raddr1_0__hier0_bF_buf5) );
BUFX4 BUFX4_39 ( .gnd(gnd), .vdd(vdd), .A(raddr1[0]), .Y(raddr1_0__hier0_bF_buf4) );
BUFX4 BUFX4_40 ( .gnd(gnd), .vdd(vdd), .A(raddr1[0]), .Y(raddr1_0__hier0_bF_buf3) );
BUFX4 BUFX4_41 ( .gnd(gnd), .vdd(vdd), .A(raddr1[0]), .Y(raddr1_0__hier0_bF_buf2) );
BUFX4 BUFX4_42 ( .gnd(gnd), .vdd(vdd), .A(raddr1[0]), .Y(raddr1_0__hier0_bF_buf1) );
BUFX4 BUFX4_43 ( .gnd(gnd), .vdd(vdd), .A(raddr1[0]), .Y(raddr1_0__hier0_bF_buf0) );
BUFX4 BUFX4_44 ( .gnd(gnd), .vdd(vdd), .A(raddr2_1_bF_buf13_), .Y(raddr2_1_bF_buf13_bF_buf3_) );
BUFX4 BUFX4_45 ( .gnd(gnd), .vdd(vdd), .A(raddr2_1_bF_buf13_), .Y(raddr2_1_bF_buf13_bF_buf2_) );
BUFX4 BUFX4_46 ( .gnd(gnd), .vdd(vdd), .A(raddr2_1_bF_buf13_), .Y(raddr2_1_bF_buf13_bF_buf1_) );
BUFX4 BUFX4_47 ( .gnd(gnd), .vdd(vdd), .A(raddr2_1_bF_buf13_), .Y(raddr2_1_bF_buf13_bF_buf0_) );
BUFX4 BUFX4_48 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf12_), .Y(raddr1_1_bF_buf12_bF_buf3_) );
BUFX4 BUFX4_49 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf12_), .Y(raddr1_1_bF_buf12_bF_buf2_) );
BUFX4 BUFX4_50 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf12_), .Y(raddr1_1_bF_buf12_bF_buf1_) );
BUFX4 BUFX4_51 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf12_), .Y(raddr1_1_bF_buf12_bF_buf0_) );
BUFX4 BUFX4_52 ( .gnd(gnd), .vdd(vdd), .A(raddr2_1_bF_buf12_), .Y(raddr2_1_bF_buf12_bF_buf3_) );
BUFX4 BUFX4_53 ( .gnd(gnd), .vdd(vdd), .A(raddr2_1_bF_buf12_), .Y(raddr2_1_bF_buf12_bF_buf2_) );
BUFX4 BUFX4_54 ( .gnd(gnd), .vdd(vdd), .A(raddr2_1_bF_buf12_), .Y(raddr2_1_bF_buf12_bF_buf1_) );
BUFX4 BUFX4_55 ( .gnd(gnd), .vdd(vdd), .A(raddr2_1_bF_buf12_), .Y(raddr2_1_bF_buf12_bF_buf0_) );
BUFX4 BUFX4_56 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf14_), .Y(raddr1_1_bF_buf14_bF_buf3_) );
BUFX4 BUFX4_57 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf14_), .Y(raddr1_1_bF_buf14_bF_buf2_) );
BUFX4 BUFX4_58 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf14_), .Y(raddr1_1_bF_buf14_bF_buf1_) );
BUFX4 BUFX4_59 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf14_), .Y(raddr1_1_bF_buf14_bF_buf0_) );
BUFX4 BUFX4_60 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf11_), .Y(raddr1_1_bF_buf11_bF_buf3_) );
BUFX4 BUFX4_61 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf11_), .Y(raddr1_1_bF_buf11_bF_buf2_) );
BUFX4 BUFX4_62 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf11_), .Y(raddr1_1_bF_buf11_bF_buf1_) );
BUFX4 BUFX4_63 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf11_), .Y(raddr1_1_bF_buf11_bF_buf0_) );
BUFX4 BUFX4_64 ( .gnd(gnd), .vdd(vdd), .A(_2101_), .Y(_2101__bF_buf7) );
BUFX4 BUFX4_65 ( .gnd(gnd), .vdd(vdd), .A(_2101_), .Y(_2101__bF_buf6) );
BUFX4 BUFX4_66 ( .gnd(gnd), .vdd(vdd), .A(_2101_), .Y(_2101__bF_buf5) );
BUFX4 BUFX4_67 ( .gnd(gnd), .vdd(vdd), .A(_2101_), .Y(_2101__bF_buf4) );
BUFX4 BUFX4_68 ( .gnd(gnd), .vdd(vdd), .A(_2101_), .Y(_2101__bF_buf3) );
BUFX4 BUFX4_69 ( .gnd(gnd), .vdd(vdd), .A(_2101_), .Y(_2101__bF_buf2) );
BUFX4 BUFX4_70 ( .gnd(gnd), .vdd(vdd), .A(_2101_), .Y(_2101__bF_buf1) );
BUFX4 BUFX4_71 ( .gnd(gnd), .vdd(vdd), .A(_2101_), .Y(_2101__bF_buf0) );
BUFX4 BUFX4_72 ( .gnd(gnd), .vdd(vdd), .A(_2365_), .Y(_2365__bF_buf4) );
BUFX4 BUFX4_73 ( .gnd(gnd), .vdd(vdd), .A(_2365_), .Y(_2365__bF_buf3) );
BUFX4 BUFX4_74 ( .gnd(gnd), .vdd(vdd), .A(_2365_), .Y(_2365__bF_buf2) );
BUFX4 BUFX4_75 ( .gnd(gnd), .vdd(vdd), .A(_2365_), .Y(_2365__bF_buf1) );
BUFX4 BUFX4_76 ( .gnd(gnd), .vdd(vdd), .A(_2365_), .Y(_2365__bF_buf0) );
BUFX4 BUFX4_77 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .Y(_1025__bF_buf3) );
BUFX4 BUFX4_78 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .Y(_1025__bF_buf2) );
BUFX4 BUFX4_79 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .Y(_1025__bF_buf1) );
BUFX4 BUFX4_80 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .Y(_1025__bF_buf0) );
BUFX4 BUFX4_81 ( .gnd(gnd), .vdd(vdd), .A(raddr2[4]), .Y(raddr2_4_bF_buf4_) );
BUFX4 BUFX4_82 ( .gnd(gnd), .vdd(vdd), .A(raddr2[4]), .Y(raddr2_4_bF_buf3_) );
BUFX4 BUFX4_83 ( .gnd(gnd), .vdd(vdd), .A(raddr2[4]), .Y(raddr2_4_bF_buf2_) );
BUFX4 BUFX4_84 ( .gnd(gnd), .vdd(vdd), .A(raddr2[4]), .Y(raddr2_4_bF_buf1_) );
BUFX4 BUFX4_85 ( .gnd(gnd), .vdd(vdd), .A(raddr2[4]), .Y(raddr2_4_bF_buf0_) );
BUFX4 BUFX4_86 ( .gnd(gnd), .vdd(vdd), .A(_1063_), .Y(_1063__bF_buf3) );
BUFX4 BUFX4_87 ( .gnd(gnd), .vdd(vdd), .A(_1063_), .Y(_1063__bF_buf2) );
BUFX4 BUFX4_88 ( .gnd(gnd), .vdd(vdd), .A(_1063_), .Y(_1063__bF_buf1) );
BUFX4 BUFX4_89 ( .gnd(gnd), .vdd(vdd), .A(_1063_), .Y(_1063__bF_buf0) );
BUFX4 BUFX4_90 ( .gnd(gnd), .vdd(vdd), .A(_1310_), .Y(_1310__bF_buf7) );
BUFX4 BUFX4_91 ( .gnd(gnd), .vdd(vdd), .A(_1310_), .Y(_1310__bF_buf6) );
BUFX4 BUFX4_92 ( .gnd(gnd), .vdd(vdd), .A(_1310_), .Y(_1310__bF_buf5) );
BUFX4 BUFX4_93 ( .gnd(gnd), .vdd(vdd), .A(_1310_), .Y(_1310__bF_buf4) );
BUFX4 BUFX4_94 ( .gnd(gnd), .vdd(vdd), .A(_1310_), .Y(_1310__bF_buf3) );
BUFX4 BUFX4_95 ( .gnd(gnd), .vdd(vdd), .A(_1310_), .Y(_1310__bF_buf2) );
BUFX4 BUFX4_96 ( .gnd(gnd), .vdd(vdd), .A(_1310_), .Y(_1310__bF_buf1) );
BUFX4 BUFX4_97 ( .gnd(gnd), .vdd(vdd), .A(_1310_), .Y(_1310__bF_buf0) );
BUFX4 BUFX4_98 ( .gnd(gnd), .vdd(vdd), .A(raddr2[1]), .Y(raddr2_1_bF_buf14_) );
BUFX4 BUFX4_99 ( .gnd(gnd), .vdd(vdd), .A(raddr2[1]), .Y(raddr2_1_bF_buf13_) );
BUFX4 BUFX4_100 ( .gnd(gnd), .vdd(vdd), .A(raddr2[1]), .Y(raddr2_1_bF_buf12_) );
BUFX4 BUFX4_101 ( .gnd(gnd), .vdd(vdd), .A(raddr2[1]), .Y(raddr2_1_bF_buf11_) );
BUFX4 BUFX4_102 ( .gnd(gnd), .vdd(vdd), .A(raddr2[1]), .Y(raddr2_1_bF_buf10_) );
BUFX4 BUFX4_103 ( .gnd(gnd), .vdd(vdd), .A(raddr2[1]), .Y(raddr2_1_bF_buf9_) );
BUFX4 BUFX4_104 ( .gnd(gnd), .vdd(vdd), .A(raddr2[1]), .Y(raddr2_1_bF_buf8_) );
BUFX4 BUFX4_105 ( .gnd(gnd), .vdd(vdd), .A(raddr2[1]), .Y(raddr2_1_bF_buf7_) );
BUFX4 BUFX4_106 ( .gnd(gnd), .vdd(vdd), .A(raddr2[1]), .Y(raddr2_1_bF_buf6_) );
BUFX4 BUFX4_107 ( .gnd(gnd), .vdd(vdd), .A(raddr2[1]), .Y(raddr2_1_bF_buf5_) );
BUFX4 BUFX4_108 ( .gnd(gnd), .vdd(vdd), .A(raddr2[1]), .Y(raddr2_1_bF_buf4_) );
BUFX4 BUFX4_109 ( .gnd(gnd), .vdd(vdd), .A(raddr2[1]), .Y(raddr2_1_bF_buf3_) );
BUFX4 BUFX4_110 ( .gnd(gnd), .vdd(vdd), .A(raddr2[1]), .Y(raddr2_1_bF_buf2_) );
BUFX4 BUFX4_111 ( .gnd(gnd), .vdd(vdd), .A(raddr2[1]), .Y(raddr2_1_bF_buf1_) );
BUFX4 BUFX4_112 ( .gnd(gnd), .vdd(vdd), .A(raddr2[1]), .Y(raddr2_1_bF_buf0_) );
BUFX4 BUFX4_113 ( .gnd(gnd), .vdd(vdd), .A(_2265_), .Y(_2265__bF_buf4) );
BUFX4 BUFX4_114 ( .gnd(gnd), .vdd(vdd), .A(_2265_), .Y(_2265__bF_buf3) );
BUFX4 BUFX4_115 ( .gnd(gnd), .vdd(vdd), .A(_2265_), .Y(_2265__bF_buf2) );
BUFX4 BUFX4_116 ( .gnd(gnd), .vdd(vdd), .A(_2265_), .Y(_2265__bF_buf1) );
BUFX4 BUFX4_117 ( .gnd(gnd), .vdd(vdd), .A(_2265_), .Y(_2265__bF_buf0) );
BUFX4 BUFX4_118 ( .gnd(gnd), .vdd(vdd), .A(raddr1[4]), .Y(raddr1_4_bF_buf4_) );
BUFX4 BUFX4_119 ( .gnd(gnd), .vdd(vdd), .A(raddr1[4]), .Y(raddr1_4_bF_buf3_) );
BUFX4 BUFX4_120 ( .gnd(gnd), .vdd(vdd), .A(raddr1[4]), .Y(raddr1_4_bF_buf2_) );
BUFX4 BUFX4_121 ( .gnd(gnd), .vdd(vdd), .A(raddr1[4]), .Y(raddr1_4_bF_buf1_) );
BUFX4 BUFX4_122 ( .gnd(gnd), .vdd(vdd), .A(raddr1[4]), .Y(raddr1_4_bF_buf0_) );
BUFX4 BUFX4_123 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .Y(_1019__bF_buf3) );
BUFX4 BUFX4_124 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .Y(_1019__bF_buf2) );
BUFX4 BUFX4_125 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .Y(_1019__bF_buf1) );
BUFX4 BUFX4_126 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .Y(_1019__bF_buf0) );
BUFX4 BUFX4_127 ( .gnd(gnd), .vdd(vdd), .A(_999_), .Y(_999__bF_buf4) );
BUFX4 BUFX4_128 ( .gnd(gnd), .vdd(vdd), .A(_999_), .Y(_999__bF_buf3) );
BUFX4 BUFX4_129 ( .gnd(gnd), .vdd(vdd), .A(_999_), .Y(_999__bF_buf2) );
BUFX4 BUFX4_130 ( .gnd(gnd), .vdd(vdd), .A(_999_), .Y(_999__bF_buf1) );
BUFX4 BUFX4_131 ( .gnd(gnd), .vdd(vdd), .A(_999_), .Y(_999__bF_buf0) );
BUFX4 BUFX4_132 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .Y(_1057__bF_buf3) );
BUFX4 BUFX4_133 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .Y(_1057__bF_buf2) );
BUFX4 BUFX4_134 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .Y(_1057__bF_buf1) );
BUFX4 BUFX4_135 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .Y(_1057__bF_buf0) );
BUFX4 BUFX4_136 ( .gnd(gnd), .vdd(vdd), .A(_2415_), .Y(_2415__bF_buf8) );
BUFX4 BUFX4_137 ( .gnd(gnd), .vdd(vdd), .A(_2415_), .Y(_2415__bF_buf7) );
BUFX4 BUFX4_138 ( .gnd(gnd), .vdd(vdd), .A(_2415_), .Y(_2415__bF_buf6) );
BUFX4 BUFX4_139 ( .gnd(gnd), .vdd(vdd), .A(_2415_), .Y(_2415__bF_buf5) );
BUFX4 BUFX4_140 ( .gnd(gnd), .vdd(vdd), .A(_2415_), .Y(_2415__bF_buf4) );
BUFX4 BUFX4_141 ( .gnd(gnd), .vdd(vdd), .A(_2415_), .Y(_2415__bF_buf3) );
BUFX4 BUFX4_142 ( .gnd(gnd), .vdd(vdd), .A(_2415_), .Y(_2415__bF_buf2) );
BUFX4 BUFX4_143 ( .gnd(gnd), .vdd(vdd), .A(_2415_), .Y(_2415__bF_buf1) );
BUFX4 BUFX4_144 ( .gnd(gnd), .vdd(vdd), .A(_2415_), .Y(_2415__bF_buf0) );
BUFX4 BUFX4_145 ( .gnd(gnd), .vdd(vdd), .A(raddr1[1]), .Y(raddr1_1_bF_buf14_) );
BUFX4 BUFX4_146 ( .gnd(gnd), .vdd(vdd), .A(raddr1[1]), .Y(raddr1_1_bF_buf13_) );
BUFX4 BUFX4_147 ( .gnd(gnd), .vdd(vdd), .A(raddr1[1]), .Y(raddr1_1_bF_buf12_) );
BUFX4 BUFX4_148 ( .gnd(gnd), .vdd(vdd), .A(raddr1[1]), .Y(raddr1_1_bF_buf11_) );
BUFX4 BUFX4_149 ( .gnd(gnd), .vdd(vdd), .A(raddr1[1]), .Y(raddr1_1_bF_buf10_) );
BUFX4 BUFX4_150 ( .gnd(gnd), .vdd(vdd), .A(raddr1[1]), .Y(raddr1_1_bF_buf9_) );
BUFX4 BUFX4_151 ( .gnd(gnd), .vdd(vdd), .A(raddr1[1]), .Y(raddr1_1_bF_buf8_) );
BUFX4 BUFX4_152 ( .gnd(gnd), .vdd(vdd), .A(raddr1[1]), .Y(raddr1_1_bF_buf7_) );
BUFX4 BUFX4_153 ( .gnd(gnd), .vdd(vdd), .A(raddr1[1]), .Y(raddr1_1_bF_buf6_) );
BUFX4 BUFX4_154 ( .gnd(gnd), .vdd(vdd), .A(raddr1[1]), .Y(raddr1_1_bF_buf5_) );
BUFX4 BUFX4_155 ( .gnd(gnd), .vdd(vdd), .A(raddr1[1]), .Y(raddr1_1_bF_buf4_) );
BUFX4 BUFX4_156 ( .gnd(gnd), .vdd(vdd), .A(raddr1[1]), .Y(raddr1_1_bF_buf3_) );
BUFX4 BUFX4_157 ( .gnd(gnd), .vdd(vdd), .A(raddr1[1]), .Y(raddr1_1_bF_buf2_) );
BUFX4 BUFX4_158 ( .gnd(gnd), .vdd(vdd), .A(raddr1[1]), .Y(raddr1_1_bF_buf1_) );
BUFX4 BUFX4_159 ( .gnd(gnd), .vdd(vdd), .A(raddr1[1]), .Y(raddr1_1_bF_buf0_) );
BUFX4 BUFX4_160 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .Y(_1571__bF_buf7) );
BUFX4 BUFX4_161 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .Y(_1571__bF_buf6) );
BUFX4 BUFX4_162 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .Y(_1571__bF_buf5) );
BUFX4 BUFX4_163 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .Y(_1571__bF_buf4) );
BUFX4 BUFX4_164 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .Y(_1571__bF_buf3) );
BUFX4 BUFX4_165 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .Y(_1571__bF_buf2) );
BUFX4 BUFX4_166 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .Y(_1571__bF_buf1) );
BUFX4 BUFX4_167 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .Y(_1571__bF_buf0) );
BUFX4 BUFX4_168 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .Y(_1207__bF_buf7) );
BUFX4 BUFX4_169 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .Y(_1207__bF_buf6) );
BUFX4 BUFX4_170 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .Y(_1207__bF_buf5) );
BUFX4 BUFX4_171 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .Y(_1207__bF_buf4) );
BUFX4 BUFX4_172 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .Y(_1207__bF_buf3) );
BUFX4 BUFX4_173 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .Y(_1207__bF_buf2) );
BUFX4 BUFX4_174 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .Y(_1207__bF_buf1) );
BUFX4 BUFX4_175 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .Y(_1207__bF_buf0) );
BUFX4 BUFX4_176 ( .gnd(gnd), .vdd(vdd), .A(_2165_), .Y(_2165__bF_buf4) );
BUFX4 BUFX4_177 ( .gnd(gnd), .vdd(vdd), .A(_2165_), .Y(_2165__bF_buf3) );
BUFX4 BUFX4_178 ( .gnd(gnd), .vdd(vdd), .A(_2165_), .Y(_2165__bF_buf2) );
BUFX4 BUFX4_179 ( .gnd(gnd), .vdd(vdd), .A(_2165_), .Y(_2165__bF_buf1) );
BUFX4 BUFX4_180 ( .gnd(gnd), .vdd(vdd), .A(_2165_), .Y(_2165__bF_buf0) );
BUFX4 BUFX4_181 ( .gnd(gnd), .vdd(vdd), .A(_1013_), .Y(_1013__bF_buf3) );
BUFX4 BUFX4_182 ( .gnd(gnd), .vdd(vdd), .A(_1013_), .Y(_1013__bF_buf2) );
BUFX4 BUFX4_183 ( .gnd(gnd), .vdd(vdd), .A(_1013_), .Y(_1013__bF_buf1) );
BUFX4 BUFX4_184 ( .gnd(gnd), .vdd(vdd), .A(_1013_), .Y(_1013__bF_buf0) );
BUFX4 BUFX4_185 ( .gnd(gnd), .vdd(vdd), .A(_1051_), .Y(_1051__bF_buf3) );
BUFX4 BUFX4_186 ( .gnd(gnd), .vdd(vdd), .A(_1051_), .Y(_1051__bF_buf2) );
BUFX4 BUFX4_187 ( .gnd(gnd), .vdd(vdd), .A(_1051_), .Y(_1051__bF_buf1) );
BUFX4 BUFX4_188 ( .gnd(gnd), .vdd(vdd), .A(_1051_), .Y(_1051__bF_buf0) );
BUFX4 BUFX4_189 ( .gnd(gnd), .vdd(vdd), .A(_1374_), .Y(_1374__bF_buf7) );
BUFX4 BUFX4_190 ( .gnd(gnd), .vdd(vdd), .A(_1374_), .Y(_1374__bF_buf6) );
BUFX4 BUFX4_191 ( .gnd(gnd), .vdd(vdd), .A(_1374_), .Y(_1374__bF_buf5) );
BUFX4 BUFX4_192 ( .gnd(gnd), .vdd(vdd), .A(_1374_), .Y(_1374__bF_buf4) );
BUFX4 BUFX4_193 ( .gnd(gnd), .vdd(vdd), .A(_1374_), .Y(_1374__bF_buf3) );
BUFX4 BUFX4_194 ( .gnd(gnd), .vdd(vdd), .A(_1374_), .Y(_1374__bF_buf2) );
BUFX4 BUFX4_195 ( .gnd(gnd), .vdd(vdd), .A(_1374_), .Y(_1374__bF_buf1) );
BUFX4 BUFX4_196 ( .gnd(gnd), .vdd(vdd), .A(_1374_), .Y(_1374__bF_buf0) );
CLKBUF1 CLKBUF1_1 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf98) );
CLKBUF1 CLKBUF1_2 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf97) );
CLKBUF1 CLKBUF1_3 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf96) );
CLKBUF1 CLKBUF1_4 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf95) );
CLKBUF1 CLKBUF1_5 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf94) );
CLKBUF1 CLKBUF1_6 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf93) );
CLKBUF1 CLKBUF1_7 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf92) );
CLKBUF1 CLKBUF1_8 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf91) );
CLKBUF1 CLKBUF1_9 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf90) );
CLKBUF1 CLKBUF1_10 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf89) );
CLKBUF1 CLKBUF1_11 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf88) );
CLKBUF1 CLKBUF1_12 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf87) );
CLKBUF1 CLKBUF1_13 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf86) );
CLKBUF1 CLKBUF1_14 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf85) );
CLKBUF1 CLKBUF1_15 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf84) );
CLKBUF1 CLKBUF1_16 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf83) );
CLKBUF1 CLKBUF1_17 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf82) );
CLKBUF1 CLKBUF1_18 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf81) );
CLKBUF1 CLKBUF1_19 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf80) );
CLKBUF1 CLKBUF1_20 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf79) );
CLKBUF1 CLKBUF1_21 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf78) );
CLKBUF1 CLKBUF1_22 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf77) );
CLKBUF1 CLKBUF1_23 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf76) );
CLKBUF1 CLKBUF1_24 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf75) );
CLKBUF1 CLKBUF1_25 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf74) );
CLKBUF1 CLKBUF1_26 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf73) );
CLKBUF1 CLKBUF1_27 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf72) );
CLKBUF1 CLKBUF1_28 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf71) );
CLKBUF1 CLKBUF1_29 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf70) );
CLKBUF1 CLKBUF1_30 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf69) );
CLKBUF1 CLKBUF1_31 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf68) );
CLKBUF1 CLKBUF1_32 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf67) );
CLKBUF1 CLKBUF1_33 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf66) );
CLKBUF1 CLKBUF1_34 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf65) );
CLKBUF1 CLKBUF1_35 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf64) );
CLKBUF1 CLKBUF1_36 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf63) );
CLKBUF1 CLKBUF1_37 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf62) );
CLKBUF1 CLKBUF1_38 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf61) );
CLKBUF1 CLKBUF1_39 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf60) );
CLKBUF1 CLKBUF1_40 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf59) );
CLKBUF1 CLKBUF1_41 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf58) );
CLKBUF1 CLKBUF1_42 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf57) );
CLKBUF1 CLKBUF1_43 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf56) );
CLKBUF1 CLKBUF1_44 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf55) );
CLKBUF1 CLKBUF1_45 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf54) );
CLKBUF1 CLKBUF1_46 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf53) );
CLKBUF1 CLKBUF1_47 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf52) );
CLKBUF1 CLKBUF1_48 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf51) );
CLKBUF1 CLKBUF1_49 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf50) );
CLKBUF1 CLKBUF1_50 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf49) );
CLKBUF1 CLKBUF1_51 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf48) );
CLKBUF1 CLKBUF1_52 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf47) );
CLKBUF1 CLKBUF1_53 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf46) );
CLKBUF1 CLKBUF1_54 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf45) );
CLKBUF1 CLKBUF1_55 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf44) );
CLKBUF1 CLKBUF1_56 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf43) );
CLKBUF1 CLKBUF1_57 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf42) );
CLKBUF1 CLKBUF1_58 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf41) );
CLKBUF1 CLKBUF1_59 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf40) );
CLKBUF1 CLKBUF1_60 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf39) );
CLKBUF1 CLKBUF1_61 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf38) );
CLKBUF1 CLKBUF1_62 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf37) );
CLKBUF1 CLKBUF1_63 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf36) );
CLKBUF1 CLKBUF1_64 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf35) );
CLKBUF1 CLKBUF1_65 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf34) );
CLKBUF1 CLKBUF1_66 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf33) );
CLKBUF1 CLKBUF1_67 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf32) );
CLKBUF1 CLKBUF1_68 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf31) );
CLKBUF1 CLKBUF1_69 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf30) );
CLKBUF1 CLKBUF1_70 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf29) );
CLKBUF1 CLKBUF1_71 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf28) );
CLKBUF1 CLKBUF1_72 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf27) );
CLKBUF1 CLKBUF1_73 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf26) );
CLKBUF1 CLKBUF1_74 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf25) );
CLKBUF1 CLKBUF1_75 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf24) );
CLKBUF1 CLKBUF1_76 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf23) );
CLKBUF1 CLKBUF1_77 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf22) );
CLKBUF1 CLKBUF1_78 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf21) );
CLKBUF1 CLKBUF1_79 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf20) );
CLKBUF1 CLKBUF1_80 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf19) );
CLKBUF1 CLKBUF1_81 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf18) );
CLKBUF1 CLKBUF1_82 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf17) );
CLKBUF1 CLKBUF1_83 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf16) );
CLKBUF1 CLKBUF1_84 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf15) );
CLKBUF1 CLKBUF1_85 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf14) );
CLKBUF1 CLKBUF1_86 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf13) );
CLKBUF1 CLKBUF1_87 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf12) );
CLKBUF1 CLKBUF1_88 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf11) );
CLKBUF1 CLKBUF1_89 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf10) );
CLKBUF1 CLKBUF1_90 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf9) );
CLKBUF1 CLKBUF1_91 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf8) );
CLKBUF1 CLKBUF1_92 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf7) );
CLKBUF1 CLKBUF1_93 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf6) );
CLKBUF1 CLKBUF1_94 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf5) );
CLKBUF1 CLKBUF1_95 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf4) );
CLKBUF1 CLKBUF1_96 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf3) );
CLKBUF1 CLKBUF1_97 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf2) );
CLKBUF1 CLKBUF1_98 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf1) );
CLKBUF1 CLKBUF1_99 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf0) );
BUFX4 BUFX4_197 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .Y(_1104__bF_buf14) );
BUFX4 BUFX4_198 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .Y(_1104__bF_buf13) );
BUFX4 BUFX4_199 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .Y(_1104__bF_buf12) );
BUFX4 BUFX4_200 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .Y(_1104__bF_buf11) );
BUFX4 BUFX4_201 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .Y(_1104__bF_buf10) );
BUFX4 BUFX4_202 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .Y(_1104__bF_buf9) );
BUFX4 BUFX4_203 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .Y(_1104__bF_buf8) );
BUFX4 BUFX4_204 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .Y(_1104__bF_buf7) );
BUFX4 BUFX4_205 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .Y(_1104__bF_buf6) );
BUFX4 BUFX4_206 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .Y(_1104__bF_buf5) );
BUFX4 BUFX4_207 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .Y(_1104__bF_buf4) );
BUFX4 BUFX4_208 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .Y(_1104__bF_buf3) );
BUFX4 BUFX4_209 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .Y(_1104__bF_buf2) );
BUFX4 BUFX4_210 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .Y(_1104__bF_buf1) );
BUFX4 BUFX4_211 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .Y(_1104__bF_buf0) );
BUFX4 BUFX4_212 ( .gnd(gnd), .vdd(vdd), .A(_1142_), .Y(_1142__bF_buf5) );
BUFX4 BUFX4_213 ( .gnd(gnd), .vdd(vdd), .A(_1142_), .Y(_1142__bF_buf4) );
BUFX4 BUFX4_214 ( .gnd(gnd), .vdd(vdd), .A(_1142_), .Y(_1142__bF_buf3) );
BUFX4 BUFX4_215 ( .gnd(gnd), .vdd(vdd), .A(_1142_), .Y(_1142__bF_buf2) );
BUFX4 BUFX4_216 ( .gnd(gnd), .vdd(vdd), .A(_1142_), .Y(_1142__bF_buf1) );
BUFX4 BUFX4_217 ( .gnd(gnd), .vdd(vdd), .A(_1142_), .Y(_1142__bF_buf0) );
BUFX4 BUFX4_218 ( .gnd(gnd), .vdd(vdd), .A(_1007_), .Y(_1007__bF_buf3) );
BUFX4 BUFX4_219 ( .gnd(gnd), .vdd(vdd), .A(_1007_), .Y(_1007__bF_buf2) );
BUFX4 BUFX4_220 ( .gnd(gnd), .vdd(vdd), .A(_1007_), .Y(_1007__bF_buf1) );
BUFX4 BUFX4_221 ( .gnd(gnd), .vdd(vdd), .A(_1007_), .Y(_1007__bF_buf0) );
BUFX4 BUFX4_222 ( .gnd(gnd), .vdd(vdd), .A(_1045_), .Y(_1045__bF_buf3) );
BUFX4 BUFX4_223 ( .gnd(gnd), .vdd(vdd), .A(_1045_), .Y(_1045__bF_buf2) );
BUFX4 BUFX4_224 ( .gnd(gnd), .vdd(vdd), .A(_1045_), .Y(_1045__bF_buf1) );
BUFX4 BUFX4_225 ( .gnd(gnd), .vdd(vdd), .A(_1045_), .Y(_1045__bF_buf0) );
BUFX4 BUFX4_226 ( .gnd(gnd), .vdd(vdd), .A(_1274_), .Y(_1274__bF_buf4) );
BUFX4 BUFX4_227 ( .gnd(gnd), .vdd(vdd), .A(_1274_), .Y(_1274__bF_buf3) );
BUFX4 BUFX4_228 ( .gnd(gnd), .vdd(vdd), .A(_1274_), .Y(_1274__bF_buf2) );
BUFX4 BUFX4_229 ( .gnd(gnd), .vdd(vdd), .A(_1274_), .Y(_1274__bF_buf1) );
BUFX4 BUFX4_230 ( .gnd(gnd), .vdd(vdd), .A(_1274_), .Y(_1274__bF_buf0) );
BUFX4 BUFX4_231 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .Y(_1039__bF_buf3) );
BUFX4 BUFX4_232 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .Y(_1039__bF_buf2) );
BUFX4 BUFX4_233 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .Y(_1039__bF_buf1) );
BUFX4 BUFX4_234 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .Y(_1039__bF_buf0) );
BUFX4 BUFX4_235 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .Y(_1803__bF_buf7) );
BUFX4 BUFX4_236 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .Y(_1803__bF_buf6) );
BUFX4 BUFX4_237 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .Y(_1803__bF_buf5) );
BUFX4 BUFX4_238 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .Y(_1803__bF_buf4) );
BUFX4 BUFX4_239 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .Y(_1803__bF_buf3) );
BUFX4 BUFX4_240 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .Y(_1803__bF_buf2) );
BUFX4 BUFX4_241 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .Y(_1803__bF_buf1) );
BUFX4 BUFX4_242 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .Y(_1803__bF_buf0) );
BUFX4 BUFX4_243 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .Y(_1001__bF_buf9) );
BUFX4 BUFX4_244 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .Y(_1001__bF_buf8) );
BUFX4 BUFX4_245 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .Y(_1001__bF_buf7) );
BUFX4 BUFX4_246 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .Y(_1001__bF_buf6) );
BUFX4 BUFX4_247 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .Y(_1001__bF_buf5) );
BUFX4 BUFX4_248 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .Y(_1001__bF_buf4) );
BUFX4 BUFX4_249 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .Y(_1001__bF_buf3) );
BUFX4 BUFX4_250 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .Y(_1001__bF_buf2) );
BUFX4 BUFX4_251 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .Y(_1001__bF_buf1) );
BUFX4 BUFX4_252 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .Y(_1001__bF_buf0) );
BUFX4 BUFX4_253 ( .gnd(gnd), .vdd(vdd), .A(_1033_), .Y(_1033__bF_buf3) );
BUFX4 BUFX4_254 ( .gnd(gnd), .vdd(vdd), .A(_1033_), .Y(_1033__bF_buf2) );
BUFX4 BUFX4_255 ( .gnd(gnd), .vdd(vdd), .A(_1033_), .Y(_1033__bF_buf1) );
BUFX4 BUFX4_256 ( .gnd(gnd), .vdd(vdd), .A(_1033_), .Y(_1033__bF_buf0) );
BUFX4 BUFX4_257 ( .gnd(gnd), .vdd(vdd), .A(_2332_), .Y(_2332__bF_buf4) );
BUFX4 BUFX4_258 ( .gnd(gnd), .vdd(vdd), .A(_2332_), .Y(_2332__bF_buf3) );
BUFX4 BUFX4_259 ( .gnd(gnd), .vdd(vdd), .A(_2332_), .Y(_2332__bF_buf2) );
BUFX4 BUFX4_260 ( .gnd(gnd), .vdd(vdd), .A(_2332_), .Y(_2332__bF_buf1) );
BUFX4 BUFX4_261 ( .gnd(gnd), .vdd(vdd), .A(_2332_), .Y(_2332__bF_buf0) );
BUFX4 BUFX4_262 ( .gnd(gnd), .vdd(vdd), .A(_1506_), .Y(_1506__bF_buf5) );
BUFX4 BUFX4_263 ( .gnd(gnd), .vdd(vdd), .A(_1506_), .Y(_1506__bF_buf4) );
BUFX4 BUFX4_264 ( .gnd(gnd), .vdd(vdd), .A(_1506_), .Y(_1506__bF_buf3) );
BUFX4 BUFX4_265 ( .gnd(gnd), .vdd(vdd), .A(_1506_), .Y(_1506__bF_buf2) );
BUFX4 BUFX4_266 ( .gnd(gnd), .vdd(vdd), .A(_1506_), .Y(_1506__bF_buf1) );
BUFX4 BUFX4_267 ( .gnd(gnd), .vdd(vdd), .A(_1506_), .Y(_1506__bF_buf0) );
BUFX4 BUFX4_268 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .Y(_1867__bF_buf4) );
BUFX4 BUFX4_269 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .Y(_1867__bF_buf3) );
BUFX4 BUFX4_270 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .Y(_1867__bF_buf2) );
BUFX4 BUFX4_271 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .Y(_1867__bF_buf1) );
BUFX4 BUFX4_272 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .Y(_1867__bF_buf0) );
BUFX4 BUFX4_273 ( .gnd(gnd), .vdd(vdd), .A(_1027_), .Y(_1027__bF_buf3) );
BUFX4 BUFX4_274 ( .gnd(gnd), .vdd(vdd), .A(_1027_), .Y(_1027__bF_buf2) );
BUFX4 BUFX4_275 ( .gnd(gnd), .vdd(vdd), .A(_1027_), .Y(_1027__bF_buf1) );
BUFX4 BUFX4_276 ( .gnd(gnd), .vdd(vdd), .A(_1027_), .Y(_1027__bF_buf0) );
BUFX4 BUFX4_277 ( .gnd(gnd), .vdd(vdd), .A(_2100_), .Y(_2100__bF_buf8) );
BUFX4 BUFX4_278 ( .gnd(gnd), .vdd(vdd), .A(_2100_), .Y(_2100__bF_buf7) );
BUFX4 BUFX4_279 ( .gnd(gnd), .vdd(vdd), .A(_2100_), .Y(_2100__bF_buf6) );
BUFX4 BUFX4_280 ( .gnd(gnd), .vdd(vdd), .A(_2100_), .Y(_2100__bF_buf5) );
BUFX4 BUFX4_281 ( .gnd(gnd), .vdd(vdd), .A(_2100_), .Y(_2100__bF_buf4) );
BUFX4 BUFX4_282 ( .gnd(gnd), .vdd(vdd), .A(_2100_), .Y(_2100__bF_buf3) );
BUFX4 BUFX4_283 ( .gnd(gnd), .vdd(vdd), .A(_2100_), .Y(_2100__bF_buf2) );
BUFX4 BUFX4_284 ( .gnd(gnd), .vdd(vdd), .A(_2100_), .Y(_2100__bF_buf1) );
BUFX4 BUFX4_285 ( .gnd(gnd), .vdd(vdd), .A(_2100_), .Y(_2100__bF_buf0) );
BUFX4 BUFX4_286 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .Y(_1309__bF_buf5) );
BUFX4 BUFX4_287 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .Y(_1309__bF_buf4) );
BUFX4 BUFX4_288 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .Y(_1309__bF_buf3) );
BUFX4 BUFX4_289 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .Y(_1309__bF_buf2) );
BUFX4 BUFX4_290 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .Y(_1309__bF_buf1) );
BUFX4 BUFX4_291 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .Y(_1309__bF_buf0) );
BUFX4 BUFX4_292 ( .gnd(gnd), .vdd(vdd), .A(_2399_), .Y(_2399__bF_buf8) );
BUFX4 BUFX4_293 ( .gnd(gnd), .vdd(vdd), .A(_2399_), .Y(_2399__bF_buf7) );
BUFX4 BUFX4_294 ( .gnd(gnd), .vdd(vdd), .A(_2399_), .Y(_2399__bF_buf6) );
BUFX4 BUFX4_295 ( .gnd(gnd), .vdd(vdd), .A(_2399_), .Y(_2399__bF_buf5) );
BUFX4 BUFX4_296 ( .gnd(gnd), .vdd(vdd), .A(_2399_), .Y(_2399__bF_buf4) );
BUFX4 BUFX4_297 ( .gnd(gnd), .vdd(vdd), .A(_2399_), .Y(_2399__bF_buf3) );
BUFX4 BUFX4_298 ( .gnd(gnd), .vdd(vdd), .A(_2399_), .Y(_2399__bF_buf2) );
BUFX4 BUFX4_299 ( .gnd(gnd), .vdd(vdd), .A(_2399_), .Y(_2399__bF_buf1) );
BUFX4 BUFX4_300 ( .gnd(gnd), .vdd(vdd), .A(_2399_), .Y(_2399__bF_buf0) );
BUFX4 BUFX4_301 ( .gnd(gnd), .vdd(vdd), .A(_1059_), .Y(_1059__bF_buf3) );
BUFX4 BUFX4_302 ( .gnd(gnd), .vdd(vdd), .A(_1059_), .Y(_1059__bF_buf2) );
BUFX4 BUFX4_303 ( .gnd(gnd), .vdd(vdd), .A(_1059_), .Y(_1059__bF_buf1) );
BUFX4 BUFX4_304 ( .gnd(gnd), .vdd(vdd), .A(_1059_), .Y(_1059__bF_buf0) );
BUFX4 BUFX4_305 ( .gnd(gnd), .vdd(vdd), .A(_2000_), .Y(_2000__bF_buf7) );
BUFX4 BUFX4_306 ( .gnd(gnd), .vdd(vdd), .A(_2000_), .Y(_2000__bF_buf6) );
BUFX4 BUFX4_307 ( .gnd(gnd), .vdd(vdd), .A(_2000_), .Y(_2000__bF_buf5) );
BUFX4 BUFX4_308 ( .gnd(gnd), .vdd(vdd), .A(_2000_), .Y(_2000__bF_buf4) );
BUFX4 BUFX4_309 ( .gnd(gnd), .vdd(vdd), .A(_2000_), .Y(_2000__bF_buf3) );
BUFX4 BUFX4_310 ( .gnd(gnd), .vdd(vdd), .A(_2000_), .Y(_2000__bF_buf2) );
BUFX4 BUFX4_311 ( .gnd(gnd), .vdd(vdd), .A(_2000_), .Y(_2000__bF_buf1) );
BUFX4 BUFX4_312 ( .gnd(gnd), .vdd(vdd), .A(_2000_), .Y(_2000__bF_buf0) );
BUFX4 BUFX4_313 ( .gnd(gnd), .vdd(vdd), .A(_1021_), .Y(_1021__bF_buf3) );
BUFX4 BUFX4_314 ( .gnd(gnd), .vdd(vdd), .A(_1021_), .Y(_1021__bF_buf2) );
BUFX4 BUFX4_315 ( .gnd(gnd), .vdd(vdd), .A(_1021_), .Y(_1021__bF_buf1) );
BUFX4 BUFX4_316 ( .gnd(gnd), .vdd(vdd), .A(_1021_), .Y(_1021__bF_buf0) );
BUFX4 BUFX4_317 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf8), .Y(raddr2_0_bF_buf96_) );
BUFX4 BUFX4_318 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf7), .Y(raddr2_0_bF_buf95_) );
BUFX4 BUFX4_319 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf6), .Y(raddr2_0_bF_buf94_) );
BUFX4 BUFX4_320 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf5), .Y(raddr2_0_bF_buf93_) );
BUFX4 BUFX4_321 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf4), .Y(raddr2_0_bF_buf92_) );
BUFX4 BUFX4_322 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf3), .Y(raddr2_0_bF_buf91_) );
BUFX4 BUFX4_323 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf2), .Y(raddr2_0_bF_buf90_) );
BUFX4 BUFX4_324 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf1), .Y(raddr2_0_bF_buf89_) );
BUFX4 BUFX4_325 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf0), .Y(raddr2_0_bF_buf88_) );
BUFX4 BUFX4_326 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf8), .Y(raddr2_0_bF_buf87_) );
BUFX4 BUFX4_327 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf7), .Y(raddr2_0_bF_buf86_) );
BUFX4 BUFX4_328 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf6), .Y(raddr2_0_bF_buf85_) );
BUFX4 BUFX4_329 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf5), .Y(raddr2_0_bF_buf84_) );
BUFX4 BUFX4_330 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf4), .Y(raddr2_0_bF_buf83_) );
BUFX4 BUFX4_331 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf3), .Y(raddr2_0_bF_buf82_) );
BUFX4 BUFX4_332 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf2), .Y(raddr2_0_bF_buf81_) );
BUFX4 BUFX4_333 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf1), .Y(raddr2_0_bF_buf80_) );
BUFX4 BUFX4_334 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf0), .Y(raddr2_0_bF_buf79_) );
BUFX4 BUFX4_335 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf8), .Y(raddr2_0_bF_buf78_) );
BUFX4 BUFX4_336 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf7), .Y(raddr2_0_bF_buf77_) );
BUFX4 BUFX4_337 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf6), .Y(raddr2_0_bF_buf76_) );
BUFX4 BUFX4_338 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf5), .Y(raddr2_0_bF_buf75_) );
BUFX4 BUFX4_339 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf4), .Y(raddr2_0_bF_buf74_) );
BUFX4 BUFX4_340 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf3), .Y(raddr2_0_bF_buf73_) );
BUFX4 BUFX4_341 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf2), .Y(raddr2_0_bF_buf72_) );
BUFX4 BUFX4_342 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf1), .Y(raddr2_0_bF_buf71_) );
BUFX4 BUFX4_343 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf0), .Y(raddr2_0_bF_buf70_) );
BUFX4 BUFX4_344 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf8), .Y(raddr2_0_bF_buf69_) );
BUFX4 BUFX4_345 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf7), .Y(raddr2_0_bF_buf68_) );
BUFX4 BUFX4_346 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf6), .Y(raddr2_0_bF_buf67_) );
BUFX4 BUFX4_347 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf5), .Y(raddr2_0_bF_buf66_) );
BUFX4 BUFX4_348 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf4), .Y(raddr2_0_bF_buf65_) );
BUFX4 BUFX4_349 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf3), .Y(raddr2_0_bF_buf64_) );
BUFX4 BUFX4_350 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf2), .Y(raddr2_0_bF_buf63_) );
BUFX4 BUFX4_351 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf1), .Y(raddr2_0_bF_buf62_) );
BUFX4 BUFX4_352 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf0), .Y(raddr2_0_bF_buf61_) );
BUFX4 BUFX4_353 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf8), .Y(raddr2_0_bF_buf60_) );
BUFX4 BUFX4_354 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf7), .Y(raddr2_0_bF_buf59_) );
BUFX4 BUFX4_355 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf6), .Y(raddr2_0_bF_buf58_) );
BUFX4 BUFX4_356 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf5), .Y(raddr2_0_bF_buf57_) );
BUFX4 BUFX4_357 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf4), .Y(raddr2_0_bF_buf56_) );
BUFX4 BUFX4_358 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf3), .Y(raddr2_0_bF_buf55_) );
BUFX4 BUFX4_359 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf2), .Y(raddr2_0_bF_buf54_) );
BUFX4 BUFX4_360 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf1), .Y(raddr2_0_bF_buf53_) );
BUFX4 BUFX4_361 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf0), .Y(raddr2_0_bF_buf52_) );
BUFX4 BUFX4_362 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf8), .Y(raddr2_0_bF_buf51_) );
BUFX4 BUFX4_363 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf7), .Y(raddr2_0_bF_buf50_) );
BUFX4 BUFX4_364 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf6), .Y(raddr2_0_bF_buf49_) );
BUFX4 BUFX4_365 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf5), .Y(raddr2_0_bF_buf48_) );
BUFX4 BUFX4_366 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf4), .Y(raddr2_0_bF_buf47_) );
BUFX4 BUFX4_367 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf3), .Y(raddr2_0_bF_buf46_) );
BUFX4 BUFX4_368 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf2), .Y(raddr2_0_bF_buf45_) );
BUFX4 BUFX4_369 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf1), .Y(raddr2_0_bF_buf44_) );
BUFX4 BUFX4_370 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf0), .Y(raddr2_0_bF_buf43_) );
BUFX4 BUFX4_371 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf8), .Y(raddr2_0_bF_buf42_) );
BUFX4 BUFX4_372 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf7), .Y(raddr2_0_bF_buf41_) );
BUFX4 BUFX4_373 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf6), .Y(raddr2_0_bF_buf40_) );
BUFX4 BUFX4_374 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf5), .Y(raddr2_0_bF_buf39_) );
BUFX4 BUFX4_375 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf4), .Y(raddr2_0_bF_buf38_) );
BUFX4 BUFX4_376 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf3), .Y(raddr2_0_bF_buf37_) );
BUFX4 BUFX4_377 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf2), .Y(raddr2_0_bF_buf36_) );
BUFX4 BUFX4_378 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf1), .Y(raddr2_0_bF_buf35_) );
BUFX4 BUFX4_379 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf0), .Y(raddr2_0_bF_buf34_) );
BUFX4 BUFX4_380 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf8), .Y(raddr2_0_bF_buf33_) );
BUFX4 BUFX4_381 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf7), .Y(raddr2_0_bF_buf32_) );
BUFX4 BUFX4_382 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf6), .Y(raddr2_0_bF_buf31_) );
BUFX4 BUFX4_383 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf5), .Y(raddr2_0_bF_buf30_) );
BUFX4 BUFX4_384 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf4), .Y(raddr2_0_bF_buf29_) );
BUFX4 BUFX4_385 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf3), .Y(raddr2_0_bF_buf28_) );
BUFX4 BUFX4_386 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf2), .Y(raddr2_0_bF_buf27_) );
BUFX4 BUFX4_387 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf1), .Y(raddr2_0_bF_buf26_) );
BUFX4 BUFX4_388 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf0), .Y(raddr2_0_bF_buf25_) );
BUFX4 BUFX4_389 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf8), .Y(raddr2_0_bF_buf24_) );
BUFX4 BUFX4_390 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf7), .Y(raddr2_0_bF_buf23_) );
BUFX4 BUFX4_391 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf6), .Y(raddr2_0_bF_buf22_) );
BUFX4 BUFX4_392 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf5), .Y(raddr2_0_bF_buf21_) );
BUFX4 BUFX4_393 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf4), .Y(raddr2_0_bF_buf20_) );
BUFX4 BUFX4_394 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf3), .Y(raddr2_0_bF_buf19_) );
BUFX4 BUFX4_395 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf2), .Y(raddr2_0_bF_buf18_) );
BUFX4 BUFX4_396 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf1), .Y(raddr2_0_bF_buf17_) );
BUFX4 BUFX4_397 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf0), .Y(raddr2_0_bF_buf16_) );
BUFX4 BUFX4_398 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf8), .Y(raddr2_0_bF_buf15_) );
BUFX4 BUFX4_399 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf7), .Y(raddr2_0_bF_buf14_) );
BUFX4 BUFX4_400 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf6), .Y(raddr2_0_bF_buf13_) );
BUFX4 BUFX4_401 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf5), .Y(raddr2_0_bF_buf12_) );
BUFX4 BUFX4_402 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf4), .Y(raddr2_0_bF_buf11_) );
BUFX4 BUFX4_403 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf3), .Y(raddr2_0_bF_buf10_) );
BUFX4 BUFX4_404 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf2), .Y(raddr2_0_bF_buf9_) );
BUFX4 BUFX4_405 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf1), .Y(raddr2_0_bF_buf8_) );
BUFX4 BUFX4_406 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf0), .Y(raddr2_0_bF_buf7_) );
BUFX4 BUFX4_407 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf8), .Y(raddr2_0_bF_buf6_) );
BUFX4 BUFX4_408 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf7), .Y(raddr2_0_bF_buf5_) );
BUFX4 BUFX4_409 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf6), .Y(raddr2_0_bF_buf4_) );
BUFX4 BUFX4_410 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf5), .Y(raddr2_0_bF_buf3_) );
BUFX4 BUFX4_411 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf4), .Y(raddr2_0_bF_buf2_) );
BUFX4 BUFX4_412 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf3), .Y(raddr2_0_bF_buf1_) );
BUFX4 BUFX4_413 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0__hier0_bF_buf2), .Y(raddr2_0_bF_buf0_) );
BUFX4 BUFX4_414 ( .gnd(gnd), .vdd(vdd), .A(_2264_), .Y(_2264__bF_buf10) );
BUFX4 BUFX4_415 ( .gnd(gnd), .vdd(vdd), .A(_2264_), .Y(_2264__bF_buf9) );
BUFX4 BUFX4_416 ( .gnd(gnd), .vdd(vdd), .A(_2264_), .Y(_2264__bF_buf8) );
BUFX4 BUFX4_417 ( .gnd(gnd), .vdd(vdd), .A(_2264_), .Y(_2264__bF_buf7) );
BUFX4 BUFX4_418 ( .gnd(gnd), .vdd(vdd), .A(_2264_), .Y(_2264__bF_buf6) );
BUFX4 BUFX4_419 ( .gnd(gnd), .vdd(vdd), .A(_2264_), .Y(_2264__bF_buf5) );
BUFX4 BUFX4_420 ( .gnd(gnd), .vdd(vdd), .A(_2264_), .Y(_2264__bF_buf4) );
BUFX4 BUFX4_421 ( .gnd(gnd), .vdd(vdd), .A(_2264_), .Y(_2264__bF_buf3) );
BUFX4 BUFX4_422 ( .gnd(gnd), .vdd(vdd), .A(_2264_), .Y(_2264__bF_buf2) );
BUFX4 BUFX4_423 ( .gnd(gnd), .vdd(vdd), .A(_2264_), .Y(_2264__bF_buf1) );
BUFX4 BUFX4_424 ( .gnd(gnd), .vdd(vdd), .A(_2264_), .Y(_2264__bF_buf0) );
BUFX4 BUFX4_425 ( .gnd(gnd), .vdd(vdd), .A(_2299_), .Y(_2299__bF_buf4) );
BUFX4 BUFX4_426 ( .gnd(gnd), .vdd(vdd), .A(_2299_), .Y(_2299__bF_buf3) );
BUFX4 BUFX4_427 ( .gnd(gnd), .vdd(vdd), .A(_2299_), .Y(_2299__bF_buf2) );
BUFX4 BUFX4_428 ( .gnd(gnd), .vdd(vdd), .A(_2299_), .Y(_2299__bF_buf1) );
BUFX4 BUFX4_429 ( .gnd(gnd), .vdd(vdd), .A(_2299_), .Y(_2299__bF_buf0) );
BUFX4 BUFX4_430 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf96_) );
BUFX4 BUFX4_431 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf95_) );
BUFX4 BUFX4_432 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf94_) );
BUFX4 BUFX4_433 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf93_) );
BUFX4 BUFX4_434 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf92_) );
BUFX4 BUFX4_435 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf91_) );
BUFX4 BUFX4_436 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf90_) );
BUFX4 BUFX4_437 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf89_) );
BUFX4 BUFX4_438 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf88_) );
BUFX4 BUFX4_439 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf87_) );
BUFX4 BUFX4_440 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf86_) );
BUFX4 BUFX4_441 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf85_) );
BUFX4 BUFX4_442 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf84_) );
BUFX4 BUFX4_443 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf83_) );
BUFX4 BUFX4_444 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf82_) );
BUFX4 BUFX4_445 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf81_) );
BUFX4 BUFX4_446 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf80_) );
BUFX4 BUFX4_447 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf79_) );
BUFX4 BUFX4_448 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf78_) );
BUFX4 BUFX4_449 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf77_) );
BUFX4 BUFX4_450 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf76_) );
BUFX4 BUFX4_451 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf75_) );
BUFX4 BUFX4_452 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf74_) );
BUFX4 BUFX4_453 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf73_) );
BUFX4 BUFX4_454 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf72_) );
BUFX4 BUFX4_455 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf71_) );
BUFX4 BUFX4_456 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf70_) );
BUFX4 BUFX4_457 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf69_) );
BUFX4 BUFX4_458 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf68_) );
BUFX4 BUFX4_459 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf67_) );
BUFX4 BUFX4_460 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf66_) );
BUFX4 BUFX4_461 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf65_) );
BUFX4 BUFX4_462 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf64_) );
BUFX4 BUFX4_463 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf63_) );
BUFX4 BUFX4_464 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf62_) );
BUFX4 BUFX4_465 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf61_) );
BUFX4 BUFX4_466 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf60_) );
BUFX4 BUFX4_467 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf59_) );
BUFX4 BUFX4_468 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf58_) );
BUFX4 BUFX4_469 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf57_) );
BUFX4 BUFX4_470 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf56_) );
BUFX4 BUFX4_471 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf55_) );
BUFX4 BUFX4_472 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf54_) );
BUFX4 BUFX4_473 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf53_) );
BUFX4 BUFX4_474 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf52_) );
BUFX4 BUFX4_475 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf51_) );
BUFX4 BUFX4_476 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf50_) );
BUFX4 BUFX4_477 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf49_) );
BUFX4 BUFX4_478 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf48_) );
BUFX4 BUFX4_479 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf47_) );
BUFX4 BUFX4_480 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf46_) );
BUFX4 BUFX4_481 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf45_) );
BUFX4 BUFX4_482 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf44_) );
BUFX4 BUFX4_483 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf43_) );
BUFX4 BUFX4_484 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf42_) );
BUFX4 BUFX4_485 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf41_) );
BUFX4 BUFX4_486 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf40_) );
BUFX4 BUFX4_487 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf39_) );
BUFX4 BUFX4_488 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf38_) );
BUFX4 BUFX4_489 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf37_) );
BUFX4 BUFX4_490 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf36_) );
BUFX4 BUFX4_491 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf35_) );
BUFX4 BUFX4_492 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf34_) );
BUFX4 BUFX4_493 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf33_) );
BUFX4 BUFX4_494 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf32_) );
BUFX4 BUFX4_495 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf31_) );
BUFX4 BUFX4_496 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf30_) );
BUFX4 BUFX4_497 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf29_) );
BUFX4 BUFX4_498 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf28_) );
BUFX4 BUFX4_499 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf27_) );
BUFX4 BUFX4_500 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf26_) );
BUFX4 BUFX4_501 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf25_) );
BUFX4 BUFX4_502 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf24_) );
BUFX4 BUFX4_503 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf23_) );
BUFX4 BUFX4_504 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf22_) );
BUFX4 BUFX4_505 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf21_) );
BUFX4 BUFX4_506 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf20_) );
BUFX4 BUFX4_507 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf19_) );
BUFX4 BUFX4_508 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf18_) );
BUFX4 BUFX4_509 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf17_) );
BUFX4 BUFX4_510 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf16_) );
BUFX4 BUFX4_511 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf15_) );
BUFX4 BUFX4_512 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf14_) );
BUFX4 BUFX4_513 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf13_) );
BUFX4 BUFX4_514 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf12_) );
BUFX4 BUFX4_515 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf11_) );
BUFX4 BUFX4_516 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf10_) );
BUFX4 BUFX4_517 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf9_) );
BUFX4 BUFX4_518 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf1), .Y(raddr1_0_bF_buf8_) );
BUFX4 BUFX4_519 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf0), .Y(raddr1_0_bF_buf7_) );
BUFX4 BUFX4_520 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf8), .Y(raddr1_0_bF_buf6_) );
BUFX4 BUFX4_521 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf7), .Y(raddr1_0_bF_buf5_) );
BUFX4 BUFX4_522 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf6), .Y(raddr1_0_bF_buf4_) );
BUFX4 BUFX4_523 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf5), .Y(raddr1_0_bF_buf3_) );
BUFX4 BUFX4_524 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf4), .Y(raddr1_0_bF_buf2_) );
BUFX4 BUFX4_525 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf3), .Y(raddr1_0_bF_buf1_) );
BUFX4 BUFX4_526 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0__hier0_bF_buf2), .Y(raddr1_0_bF_buf0_) );
BUFX4 BUFX4_527 ( .gnd(gnd), .vdd(vdd), .A(_1015_), .Y(_1015__bF_buf3) );
BUFX4 BUFX4_528 ( .gnd(gnd), .vdd(vdd), .A(_1015_), .Y(_1015__bF_buf2) );
BUFX4 BUFX4_529 ( .gnd(gnd), .vdd(vdd), .A(_1015_), .Y(_1015__bF_buf1) );
BUFX4 BUFX4_530 ( .gnd(gnd), .vdd(vdd), .A(_1015_), .Y(_1015__bF_buf0) );
BUFX4 BUFX4_531 ( .gnd(gnd), .vdd(vdd), .A(_1053_), .Y(_1053__bF_buf3) );
BUFX4 BUFX4_532 ( .gnd(gnd), .vdd(vdd), .A(_1053_), .Y(_1053__bF_buf2) );
BUFX4 BUFX4_533 ( .gnd(gnd), .vdd(vdd), .A(_1053_), .Y(_1053__bF_buf1) );
BUFX4 BUFX4_534 ( .gnd(gnd), .vdd(vdd), .A(_1053_), .Y(_1053__bF_buf0) );
BUFX4 BUFX4_535 ( .gnd(gnd), .vdd(vdd), .A(_992_), .Y(_992__bF_buf3) );
BUFX4 BUFX4_536 ( .gnd(gnd), .vdd(vdd), .A(_992_), .Y(_992__bF_buf2) );
BUFX4 BUFX4_537 ( .gnd(gnd), .vdd(vdd), .A(_992_), .Y(_992__bF_buf1) );
BUFX4 BUFX4_538 ( .gnd(gnd), .vdd(vdd), .A(_992_), .Y(_992__bF_buf0) );
BUFX4 BUFX4_539 ( .gnd(gnd), .vdd(vdd), .A(_2064_), .Y(_2064__bF_buf4) );
BUFX4 BUFX4_540 ( .gnd(gnd), .vdd(vdd), .A(_2064_), .Y(_2064__bF_buf3) );
BUFX4 BUFX4_541 ( .gnd(gnd), .vdd(vdd), .A(_2064_), .Y(_2064__bF_buf2) );
BUFX4 BUFX4_542 ( .gnd(gnd), .vdd(vdd), .A(_2064_), .Y(_2064__bF_buf1) );
BUFX4 BUFX4_543 ( .gnd(gnd), .vdd(vdd), .A(_2064_), .Y(_2064__bF_buf0) );
BUFX4 BUFX4_544 ( .gnd(gnd), .vdd(vdd), .A(_1009_), .Y(_1009__bF_buf3) );
BUFX4 BUFX4_545 ( .gnd(gnd), .vdd(vdd), .A(_1009_), .Y(_1009__bF_buf2) );
BUFX4 BUFX4_546 ( .gnd(gnd), .vdd(vdd), .A(_1009_), .Y(_1009__bF_buf1) );
BUFX4 BUFX4_547 ( .gnd(gnd), .vdd(vdd), .A(_1009_), .Y(_1009__bF_buf0) );
BUFX4 BUFX4_548 ( .gnd(gnd), .vdd(vdd), .A(_1047_), .Y(_1047__bF_buf3) );
BUFX4 BUFX4_549 ( .gnd(gnd), .vdd(vdd), .A(_1047_), .Y(_1047__bF_buf2) );
BUFX4 BUFX4_550 ( .gnd(gnd), .vdd(vdd), .A(_1047_), .Y(_1047__bF_buf1) );
BUFX4 BUFX4_551 ( .gnd(gnd), .vdd(vdd), .A(_1047_), .Y(_1047__bF_buf0) );
BUFX4 BUFX4_552 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .Y(_1141__bF_buf7) );
BUFX4 BUFX4_553 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .Y(_1141__bF_buf6) );
BUFX4 BUFX4_554 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .Y(_1141__bF_buf5) );
BUFX4 BUFX4_555 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .Y(_1141__bF_buf4) );
BUFX4 BUFX4_556 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .Y(_1141__bF_buf3) );
BUFX4 BUFX4_557 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .Y(_1141__bF_buf2) );
BUFX4 BUFX4_558 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .Y(_1141__bF_buf1) );
BUFX4 BUFX4_559 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .Y(_1141__bF_buf0) );
BUFX4 BUFX4_560 ( .gnd(gnd), .vdd(vdd), .A(_1902_), .Y(_1902__bF_buf7) );
BUFX4 BUFX4_561 ( .gnd(gnd), .vdd(vdd), .A(_1902_), .Y(_1902__bF_buf6) );
BUFX4 BUFX4_562 ( .gnd(gnd), .vdd(vdd), .A(_1902_), .Y(_1902__bF_buf5) );
BUFX4 BUFX4_563 ( .gnd(gnd), .vdd(vdd), .A(_1902_), .Y(_1902__bF_buf4) );
BUFX4 BUFX4_564 ( .gnd(gnd), .vdd(vdd), .A(_1902_), .Y(_1902__bF_buf3) );
BUFX4 BUFX4_565 ( .gnd(gnd), .vdd(vdd), .A(_1902_), .Y(_1902__bF_buf2) );
BUFX4 BUFX4_566 ( .gnd(gnd), .vdd(vdd), .A(_1902_), .Y(_1902__bF_buf1) );
BUFX4 BUFX4_567 ( .gnd(gnd), .vdd(vdd), .A(_1902_), .Y(_1902__bF_buf0) );
BUFX4 BUFX4_568 ( .gnd(gnd), .vdd(vdd), .A(_1003_), .Y(_1003__bF_buf3) );
BUFX4 BUFX4_569 ( .gnd(gnd), .vdd(vdd), .A(_1003_), .Y(_1003__bF_buf2) );
BUFX4 BUFX4_570 ( .gnd(gnd), .vdd(vdd), .A(_1003_), .Y(_1003__bF_buf1) );
BUFX4 BUFX4_571 ( .gnd(gnd), .vdd(vdd), .A(_1003_), .Y(_1003__bF_buf0) );
BUFX4 BUFX4_572 ( .gnd(gnd), .vdd(vdd), .A(_1041_), .Y(_1041__bF_buf3) );
BUFX4 BUFX4_573 ( .gnd(gnd), .vdd(vdd), .A(_1041_), .Y(_1041__bF_buf2) );
BUFX4 BUFX4_574 ( .gnd(gnd), .vdd(vdd), .A(_1041_), .Y(_1041__bF_buf1) );
BUFX4 BUFX4_575 ( .gnd(gnd), .vdd(vdd), .A(_1041_), .Y(_1041__bF_buf0) );
BUFX4 BUFX4_576 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf7) );
BUFX4 BUFX4_577 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf6) );
BUFX4 BUFX4_578 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf5) );
BUFX4 BUFX4_579 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf4) );
BUFX4 BUFX4_580 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf3) );
BUFX4 BUFX4_581 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf2) );
BUFX4 BUFX4_582 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf1) );
BUFX4 BUFX4_583 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .Y(_1000__bF_buf0) );
BUFX4 BUFX4_584 ( .gnd(gnd), .vdd(vdd), .A(_1705_), .Y(_1705__bF_buf7) );
BUFX4 BUFX4_585 ( .gnd(gnd), .vdd(vdd), .A(_1705_), .Y(_1705__bF_buf6) );
BUFX4 BUFX4_586 ( .gnd(gnd), .vdd(vdd), .A(_1705_), .Y(_1705__bF_buf5) );
BUFX4 BUFX4_587 ( .gnd(gnd), .vdd(vdd), .A(_1705_), .Y(_1705__bF_buf4) );
BUFX4 BUFX4_588 ( .gnd(gnd), .vdd(vdd), .A(_1705_), .Y(_1705__bF_buf3) );
BUFX4 BUFX4_589 ( .gnd(gnd), .vdd(vdd), .A(_1705_), .Y(_1705__bF_buf2) );
BUFX4 BUFX4_590 ( .gnd(gnd), .vdd(vdd), .A(_1705_), .Y(_1705__bF_buf1) );
BUFX4 BUFX4_591 ( .gnd(gnd), .vdd(vdd), .A(_1705_), .Y(_1705__bF_buf0) );
BUFX4 BUFX4_592 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .Y(_1035__bF_buf3) );
BUFX4 BUFX4_593 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .Y(_1035__bF_buf2) );
BUFX4 BUFX4_594 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .Y(_1035__bF_buf1) );
BUFX4 BUFX4_595 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .Y(_1035__bF_buf0) );
BUFX4 BUFX4_596 ( .gnd(gnd), .vdd(vdd), .A(_1605_), .Y(_1605__bF_buf7) );
BUFX4 BUFX4_597 ( .gnd(gnd), .vdd(vdd), .A(_1605_), .Y(_1605__bF_buf6) );
BUFX4 BUFX4_598 ( .gnd(gnd), .vdd(vdd), .A(_1605_), .Y(_1605__bF_buf5) );
BUFX4 BUFX4_599 ( .gnd(gnd), .vdd(vdd), .A(_1605_), .Y(_1605__bF_buf4) );
BUFX4 BUFX4_600 ( .gnd(gnd), .vdd(vdd), .A(_1605_), .Y(_1605__bF_buf3) );
BUFX4 BUFX4_601 ( .gnd(gnd), .vdd(vdd), .A(_1605_), .Y(_1605__bF_buf2) );
BUFX4 BUFX4_602 ( .gnd(gnd), .vdd(vdd), .A(_1605_), .Y(_1605__bF_buf1) );
BUFX4 BUFX4_603 ( .gnd(gnd), .vdd(vdd), .A(_1605_), .Y(_1605__bF_buf0) );
BUFX4 BUFX4_604 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .Y(_1070__bF_buf10) );
BUFX4 BUFX4_605 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .Y(_1070__bF_buf9) );
BUFX4 BUFX4_606 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .Y(_1070__bF_buf8) );
BUFX4 BUFX4_607 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .Y(_1070__bF_buf7) );
BUFX4 BUFX4_608 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .Y(_1070__bF_buf6) );
BUFX4 BUFX4_609 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .Y(_1070__bF_buf5) );
BUFX4 BUFX4_610 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .Y(_1070__bF_buf4) );
BUFX4 BUFX4_611 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .Y(_1070__bF_buf3) );
BUFX4 BUFX4_612 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .Y(_1070__bF_buf2) );
BUFX4 BUFX4_613 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .Y(_1070__bF_buf1) );
BUFX4 BUFX4_614 ( .gnd(gnd), .vdd(vdd), .A(_1070_), .Y(_1070__bF_buf0) );
BUFX4 BUFX4_615 ( .gnd(gnd), .vdd(vdd), .A(_1966_), .Y(_1966__bF_buf7) );
BUFX4 BUFX4_616 ( .gnd(gnd), .vdd(vdd), .A(_1966_), .Y(_1966__bF_buf6) );
BUFX4 BUFX4_617 ( .gnd(gnd), .vdd(vdd), .A(_1966_), .Y(_1966__bF_buf5) );
BUFX4 BUFX4_618 ( .gnd(gnd), .vdd(vdd), .A(_1966_), .Y(_1966__bF_buf4) );
BUFX4 BUFX4_619 ( .gnd(gnd), .vdd(vdd), .A(_1966_), .Y(_1966__bF_buf3) );
BUFX4 BUFX4_620 ( .gnd(gnd), .vdd(vdd), .A(_1966_), .Y(_1966__bF_buf2) );
BUFX4 BUFX4_621 ( .gnd(gnd), .vdd(vdd), .A(_1966_), .Y(_1966__bF_buf1) );
BUFX4 BUFX4_622 ( .gnd(gnd), .vdd(vdd), .A(_1966_), .Y(_1966__bF_buf0) );
BUFX4 BUFX4_623 ( .gnd(gnd), .vdd(vdd), .A(_1029_), .Y(_1029__bF_buf3) );
BUFX4 BUFX4_624 ( .gnd(gnd), .vdd(vdd), .A(_1029_), .Y(_1029__bF_buf2) );
BUFX4 BUFX4_625 ( .gnd(gnd), .vdd(vdd), .A(_1029_), .Y(_1029__bF_buf1) );
BUFX4 BUFX4_626 ( .gnd(gnd), .vdd(vdd), .A(_1029_), .Y(_1029__bF_buf0) );
BUFX4 BUFX4_627 ( .gnd(gnd), .vdd(vdd), .A(_4036_), .Y(_4036__bF_buf8) );
BUFX4 BUFX4_628 ( .gnd(gnd), .vdd(vdd), .A(_4036_), .Y(_4036__bF_buf7) );
BUFX4 BUFX4_629 ( .gnd(gnd), .vdd(vdd), .A(_4036_), .Y(_4036__bF_buf6) );
BUFX4 BUFX4_630 ( .gnd(gnd), .vdd(vdd), .A(_4036_), .Y(_4036__bF_buf5) );
BUFX4 BUFX4_631 ( .gnd(gnd), .vdd(vdd), .A(_4036_), .Y(_4036__bF_buf4) );
BUFX4 BUFX4_632 ( .gnd(gnd), .vdd(vdd), .A(_4036_), .Y(_4036__bF_buf3) );
BUFX4 BUFX4_633 ( .gnd(gnd), .vdd(vdd), .A(_4036_), .Y(_4036__bF_buf2) );
BUFX4 BUFX4_634 ( .gnd(gnd), .vdd(vdd), .A(_4036_), .Y(_4036__bF_buf1) );
BUFX4 BUFX4_635 ( .gnd(gnd), .vdd(vdd), .A(_4036_), .Y(_4036__bF_buf0) );
BUFX4 BUFX4_636 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .Y(_1408__bF_buf7) );
BUFX4 BUFX4_637 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .Y(_1408__bF_buf6) );
BUFX4 BUFX4_638 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .Y(_1408__bF_buf5) );
BUFX4 BUFX4_639 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .Y(_1408__bF_buf4) );
BUFX4 BUFX4_640 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .Y(_1408__bF_buf3) );
BUFX4 BUFX4_641 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .Y(_1408__bF_buf2) );
BUFX4 BUFX4_642 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .Y(_1408__bF_buf1) );
BUFX4 BUFX4_643 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .Y(_1408__bF_buf0) );
BUFX4 BUFX4_644 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .Y(_1769__bF_buf7) );
BUFX4 BUFX4_645 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .Y(_1769__bF_buf6) );
BUFX4 BUFX4_646 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .Y(_1769__bF_buf5) );
BUFX4 BUFX4_647 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .Y(_1769__bF_buf4) );
BUFX4 BUFX4_648 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .Y(_1769__bF_buf3) );
BUFX4 BUFX4_649 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .Y(_1769__bF_buf2) );
BUFX4 BUFX4_650 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .Y(_1769__bF_buf1) );
BUFX4 BUFX4_651 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .Y(_1769__bF_buf0) );
BUFX4 BUFX4_652 ( .gnd(gnd), .vdd(vdd), .A(_4033_), .Y(_4033__bF_buf7) );
BUFX4 BUFX4_653 ( .gnd(gnd), .vdd(vdd), .A(_4033_), .Y(_4033__bF_buf6) );
BUFX4 BUFX4_654 ( .gnd(gnd), .vdd(vdd), .A(_4033_), .Y(_4033__bF_buf5) );
BUFX4 BUFX4_655 ( .gnd(gnd), .vdd(vdd), .A(_4033_), .Y(_4033__bF_buf4) );
BUFX4 BUFX4_656 ( .gnd(gnd), .vdd(vdd), .A(_4033_), .Y(_4033__bF_buf3) );
BUFX4 BUFX4_657 ( .gnd(gnd), .vdd(vdd), .A(_4033_), .Y(_4033__bF_buf2) );
BUFX4 BUFX4_658 ( .gnd(gnd), .vdd(vdd), .A(_4033_), .Y(_4033__bF_buf1) );
BUFX4 BUFX4_659 ( .gnd(gnd), .vdd(vdd), .A(_4033_), .Y(_4033__bF_buf0) );
BUFX4 BUFX4_660 ( .gnd(gnd), .vdd(vdd), .A(_2231_), .Y(_2231__bF_buf4) );
BUFX4 BUFX4_661 ( .gnd(gnd), .vdd(vdd), .A(_2231_), .Y(_2231__bF_buf3) );
BUFX4 BUFX4_662 ( .gnd(gnd), .vdd(vdd), .A(_2231_), .Y(_2231__bF_buf2) );
BUFX4 BUFX4_663 ( .gnd(gnd), .vdd(vdd), .A(_2231_), .Y(_2231__bF_buf1) );
BUFX4 BUFX4_664 ( .gnd(gnd), .vdd(vdd), .A(_2231_), .Y(_2231__bF_buf0) );
BUFX4 BUFX4_665 ( .gnd(gnd), .vdd(vdd), .A(_1023_), .Y(_1023__bF_buf3) );
BUFX4 BUFX4_666 ( .gnd(gnd), .vdd(vdd), .A(_1023_), .Y(_1023__bF_buf2) );
BUFX4 BUFX4_667 ( .gnd(gnd), .vdd(vdd), .A(_1023_), .Y(_1023__bF_buf1) );
BUFX4 BUFX4_668 ( .gnd(gnd), .vdd(vdd), .A(_1023_), .Y(_1023__bF_buf0) );
BUFX4 BUFX4_669 ( .gnd(gnd), .vdd(vdd), .A(raddr2[2]), .Y(raddr2_2_bF_buf10_) );
BUFX4 BUFX4_670 ( .gnd(gnd), .vdd(vdd), .A(raddr2[2]), .Y(raddr2_2_bF_buf9_) );
BUFX4 BUFX4_671 ( .gnd(gnd), .vdd(vdd), .A(raddr2[2]), .Y(raddr2_2_bF_buf8_) );
BUFX4 BUFX4_672 ( .gnd(gnd), .vdd(vdd), .A(raddr2[2]), .Y(raddr2_2_bF_buf7_) );
BUFX4 BUFX4_673 ( .gnd(gnd), .vdd(vdd), .A(raddr2[2]), .Y(raddr2_2_bF_buf6_) );
BUFX4 BUFX4_674 ( .gnd(gnd), .vdd(vdd), .A(raddr2[2]), .Y(raddr2_2_bF_buf5_) );
BUFX4 BUFX4_675 ( .gnd(gnd), .vdd(vdd), .A(raddr2[2]), .Y(raddr2_2_bF_buf4_) );
BUFX4 BUFX4_676 ( .gnd(gnd), .vdd(vdd), .A(raddr2[2]), .Y(raddr2_2_bF_buf3_) );
BUFX4 BUFX4_677 ( .gnd(gnd), .vdd(vdd), .A(raddr2[2]), .Y(raddr2_2_bF_buf2_) );
BUFX4 BUFX4_678 ( .gnd(gnd), .vdd(vdd), .A(raddr2[2]), .Y(raddr2_2_bF_buf1_) );
BUFX4 BUFX4_679 ( .gnd(gnd), .vdd(vdd), .A(raddr2[2]), .Y(raddr2_2_bF_buf0_) );
BUFX4 BUFX4_680 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .Y(_1061__bF_buf3) );
BUFX4 BUFX4_681 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .Y(_1061__bF_buf2) );
BUFX4 BUFX4_682 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .Y(_1061__bF_buf1) );
BUFX4 BUFX4_683 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .Y(_1061__bF_buf0) );
BUFX4 BUFX4_684 ( .gnd(gnd), .vdd(vdd), .A(_2398_), .Y(_2398__bF_buf7) );
BUFX4 BUFX4_685 ( .gnd(gnd), .vdd(vdd), .A(_2398_), .Y(_2398__bF_buf6) );
BUFX4 BUFX4_686 ( .gnd(gnd), .vdd(vdd), .A(_2398_), .Y(_2398__bF_buf5) );
BUFX4 BUFX4_687 ( .gnd(gnd), .vdd(vdd), .A(_2398_), .Y(_2398__bF_buf4) );
BUFX4 BUFX4_688 ( .gnd(gnd), .vdd(vdd), .A(_2398_), .Y(_2398__bF_buf3) );
BUFX4 BUFX4_689 ( .gnd(gnd), .vdd(vdd), .A(_2398_), .Y(_2398__bF_buf2) );
BUFX4 BUFX4_690 ( .gnd(gnd), .vdd(vdd), .A(_2398_), .Y(_2398__bF_buf1) );
BUFX4 BUFX4_691 ( .gnd(gnd), .vdd(vdd), .A(_2398_), .Y(_2398__bF_buf0) );
BUFX4 BUFX4_692 ( .gnd(gnd), .vdd(vdd), .A(_1669_), .Y(_1669__bF_buf4) );
BUFX4 BUFX4_693 ( .gnd(gnd), .vdd(vdd), .A(_1669_), .Y(_1669__bF_buf3) );
BUFX4 BUFX4_694 ( .gnd(gnd), .vdd(vdd), .A(_1669_), .Y(_1669__bF_buf2) );
BUFX4 BUFX4_695 ( .gnd(gnd), .vdd(vdd), .A(_1669_), .Y(_1669__bF_buf1) );
BUFX4 BUFX4_696 ( .gnd(gnd), .vdd(vdd), .A(_1669_), .Y(_1669__bF_buf0) );
BUFX4 BUFX4_697 ( .gnd(gnd), .vdd(vdd), .A(raddr1[2]), .Y(raddr1_2_bF_buf10_) );
BUFX4 BUFX4_698 ( .gnd(gnd), .vdd(vdd), .A(raddr1[2]), .Y(raddr1_2_bF_buf9_) );
BUFX4 BUFX4_699 ( .gnd(gnd), .vdd(vdd), .A(raddr1[2]), .Y(raddr1_2_bF_buf8_) );
BUFX4 BUFX4_700 ( .gnd(gnd), .vdd(vdd), .A(raddr1[2]), .Y(raddr1_2_bF_buf7_) );
BUFX4 BUFX4_701 ( .gnd(gnd), .vdd(vdd), .A(raddr1[2]), .Y(raddr1_2_bF_buf6_) );
BUFX4 BUFX4_702 ( .gnd(gnd), .vdd(vdd), .A(raddr1[2]), .Y(raddr1_2_bF_buf5_) );
BUFX4 BUFX4_703 ( .gnd(gnd), .vdd(vdd), .A(raddr1[2]), .Y(raddr1_2_bF_buf4_) );
BUFX4 BUFX4_704 ( .gnd(gnd), .vdd(vdd), .A(raddr1[2]), .Y(raddr1_2_bF_buf3_) );
BUFX4 BUFX4_705 ( .gnd(gnd), .vdd(vdd), .A(raddr1[2]), .Y(raddr1_2_bF_buf2_) );
BUFX4 BUFX4_706 ( .gnd(gnd), .vdd(vdd), .A(raddr1[2]), .Y(raddr1_2_bF_buf1_) );
BUFX4 BUFX4_707 ( .gnd(gnd), .vdd(vdd), .A(raddr1[2]), .Y(raddr1_2_bF_buf0_) );
BUFX4 BUFX4_708 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .Y(_1017__bF_buf3) );
BUFX4 BUFX4_709 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .Y(_1017__bF_buf2) );
BUFX4 BUFX4_710 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .Y(_1017__bF_buf1) );
BUFX4 BUFX4_711 ( .gnd(gnd), .vdd(vdd), .A(_1017_), .Y(_1017__bF_buf0) );
BUFX4 BUFX4_712 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .Y(_1055__bF_buf3) );
BUFX4 BUFX4_713 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .Y(_1055__bF_buf2) );
BUFX4 BUFX4_714 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .Y(_1055__bF_buf1) );
BUFX4 BUFX4_715 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .Y(_1055__bF_buf0) );
BUFX4 BUFX4_716 ( .gnd(gnd), .vdd(vdd), .A(_1472_), .Y(_1472__bF_buf4) );
BUFX4 BUFX4_717 ( .gnd(gnd), .vdd(vdd), .A(_1472_), .Y(_1472__bF_buf3) );
BUFX4 BUFX4_718 ( .gnd(gnd), .vdd(vdd), .A(_1472_), .Y(_1472__bF_buf2) );
BUFX4 BUFX4_719 ( .gnd(gnd), .vdd(vdd), .A(_1472_), .Y(_1472__bF_buf1) );
BUFX4 BUFX4_720 ( .gnd(gnd), .vdd(vdd), .A(_1472_), .Y(_1472__bF_buf0) );
BUFX4 BUFX4_721 ( .gnd(gnd), .vdd(vdd), .A(_2198_), .Y(_2198__bF_buf4) );
BUFX4 BUFX4_722 ( .gnd(gnd), .vdd(vdd), .A(_2198_), .Y(_2198__bF_buf3) );
BUFX4 BUFX4_723 ( .gnd(gnd), .vdd(vdd), .A(_2198_), .Y(_2198__bF_buf2) );
BUFX4 BUFX4_724 ( .gnd(gnd), .vdd(vdd), .A(_2198_), .Y(_2198__bF_buf1) );
BUFX4 BUFX4_725 ( .gnd(gnd), .vdd(vdd), .A(_2198_), .Y(_2198__bF_buf0) );
BUFX4 BUFX4_726 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .Y(_1049__bF_buf3) );
BUFX4 BUFX4_727 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .Y(_1049__bF_buf2) );
BUFX4 BUFX4_728 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .Y(_1049__bF_buf1) );
BUFX4 BUFX4_729 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .Y(_1049__bF_buf0) );
BUFX4 BUFX4_730 ( .gnd(gnd), .vdd(vdd), .A(_1011_), .Y(_1011__bF_buf3) );
BUFX4 BUFX4_731 ( .gnd(gnd), .vdd(vdd), .A(_1011_), .Y(_1011__bF_buf2) );
BUFX4 BUFX4_732 ( .gnd(gnd), .vdd(vdd), .A(_1011_), .Y(_1011__bF_buf1) );
BUFX4 BUFX4_733 ( .gnd(gnd), .vdd(vdd), .A(_1011_), .Y(_1011__bF_buf0) );
BUFX4 BUFX4_734 ( .gnd(gnd), .vdd(vdd), .A(_1240_), .Y(_1240__bF_buf4) );
BUFX4 BUFX4_735 ( .gnd(gnd), .vdd(vdd), .A(_1240_), .Y(_1240__bF_buf3) );
BUFX4 BUFX4_736 ( .gnd(gnd), .vdd(vdd), .A(_1240_), .Y(_1240__bF_buf2) );
BUFX4 BUFX4_737 ( .gnd(gnd), .vdd(vdd), .A(_1240_), .Y(_1240__bF_buf1) );
BUFX4 BUFX4_738 ( .gnd(gnd), .vdd(vdd), .A(_1240_), .Y(_1240__bF_buf0) );
BUFX4 BUFX4_739 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .Y(_1105__bF_buf7) );
BUFX4 BUFX4_740 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .Y(_1105__bF_buf6) );
BUFX4 BUFX4_741 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .Y(_1105__bF_buf5) );
BUFX4 BUFX4_742 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .Y(_1105__bF_buf4) );
BUFX4 BUFX4_743 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .Y(_1105__bF_buf3) );
BUFX4 BUFX4_744 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .Y(_1105__bF_buf2) );
BUFX4 BUFX4_745 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .Y(_1105__bF_buf1) );
BUFX4 BUFX4_746 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .Y(_1105__bF_buf0) );
BUFX4 BUFX4_747 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .Y(_1143__bF_buf7) );
BUFX4 BUFX4_748 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .Y(_1143__bF_buf6) );
BUFX4 BUFX4_749 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .Y(_1143__bF_buf5) );
BUFX4 BUFX4_750 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .Y(_1143__bF_buf4) );
BUFX4 BUFX4_751 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .Y(_1143__bF_buf3) );
BUFX4 BUFX4_752 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .Y(_1143__bF_buf2) );
BUFX4 BUFX4_753 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .Y(_1143__bF_buf1) );
BUFX4 BUFX4_754 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .Y(_1143__bF_buf0) );
BUFX4 BUFX4_755 ( .gnd(gnd), .vdd(vdd), .A(_1005_), .Y(_1005__bF_buf3) );
BUFX4 BUFX4_756 ( .gnd(gnd), .vdd(vdd), .A(_1005_), .Y(_1005__bF_buf2) );
BUFX4 BUFX4_757 ( .gnd(gnd), .vdd(vdd), .A(_1005_), .Y(_1005__bF_buf1) );
BUFX4 BUFX4_758 ( .gnd(gnd), .vdd(vdd), .A(_1005_), .Y(_1005__bF_buf0) );
BUFX4 BUFX4_759 ( .gnd(gnd), .vdd(vdd), .A(_1043_), .Y(_1043__bF_buf3) );
BUFX4 BUFX4_760 ( .gnd(gnd), .vdd(vdd), .A(_1043_), .Y(_1043__bF_buf2) );
BUFX4 BUFX4_761 ( .gnd(gnd), .vdd(vdd), .A(_1043_), .Y(_1043__bF_buf1) );
BUFX4 BUFX4_762 ( .gnd(gnd), .vdd(vdd), .A(_1043_), .Y(_1043__bF_buf0) );
BUFX4 BUFX4_763 ( .gnd(gnd), .vdd(vdd), .A(_1901_), .Y(_1901__bF_buf5) );
BUFX4 BUFX4_764 ( .gnd(gnd), .vdd(vdd), .A(_1901_), .Y(_1901__bF_buf4) );
BUFX4 BUFX4_765 ( .gnd(gnd), .vdd(vdd), .A(_1901_), .Y(_1901__bF_buf3) );
BUFX4 BUFX4_766 ( .gnd(gnd), .vdd(vdd), .A(_1901_), .Y(_1901__bF_buf2) );
BUFX4 BUFX4_767 ( .gnd(gnd), .vdd(vdd), .A(_1901_), .Y(_1901__bF_buf1) );
BUFX4 BUFX4_768 ( .gnd(gnd), .vdd(vdd), .A(_1901_), .Y(_1901__bF_buf0) );
BUFX4 BUFX4_769 ( .gnd(gnd), .vdd(vdd), .A(_1037_), .Y(_1037__bF_buf3) );
BUFX4 BUFX4_770 ( .gnd(gnd), .vdd(vdd), .A(_1037_), .Y(_1037__bF_buf2) );
BUFX4 BUFX4_771 ( .gnd(gnd), .vdd(vdd), .A(_1037_), .Y(_1037__bF_buf1) );
BUFX4 BUFX4_772 ( .gnd(gnd), .vdd(vdd), .A(_1037_), .Y(_1037__bF_buf0) );
BUFX4 BUFX4_773 ( .gnd(gnd), .vdd(vdd), .A(_1704_), .Y(_1704__bF_buf5) );
BUFX4 BUFX4_774 ( .gnd(gnd), .vdd(vdd), .A(_1704_), .Y(_1704__bF_buf4) );
BUFX4 BUFX4_775 ( .gnd(gnd), .vdd(vdd), .A(_1704_), .Y(_1704__bF_buf3) );
BUFX4 BUFX4_776 ( .gnd(gnd), .vdd(vdd), .A(_1704_), .Y(_1704__bF_buf2) );
BUFX4 BUFX4_777 ( .gnd(gnd), .vdd(vdd), .A(_1704_), .Y(_1704__bF_buf1) );
BUFX4 BUFX4_778 ( .gnd(gnd), .vdd(vdd), .A(_1704_), .Y(_1704__bF_buf0) );
BUFX4 BUFX4_779 ( .gnd(gnd), .vdd(vdd), .A(_1069_), .Y(_1069__bF_buf4) );
BUFX4 BUFX4_780 ( .gnd(gnd), .vdd(vdd), .A(_1069_), .Y(_1069__bF_buf3) );
BUFX4 BUFX4_781 ( .gnd(gnd), .vdd(vdd), .A(_1069_), .Y(_1069__bF_buf2) );
BUFX4 BUFX4_782 ( .gnd(gnd), .vdd(vdd), .A(_1069_), .Y(_1069__bF_buf1) );
BUFX4 BUFX4_783 ( .gnd(gnd), .vdd(vdd), .A(_1069_), .Y(_1069__bF_buf0) );
BUFX4 BUFX4_784 ( .gnd(gnd), .vdd(vdd), .A(_4038_), .Y(_4038__bF_buf8) );
BUFX4 BUFX4_785 ( .gnd(gnd), .vdd(vdd), .A(_4038_), .Y(_4038__bF_buf7) );
BUFX4 BUFX4_786 ( .gnd(gnd), .vdd(vdd), .A(_4038_), .Y(_4038__bF_buf6) );
BUFX4 BUFX4_787 ( .gnd(gnd), .vdd(vdd), .A(_4038_), .Y(_4038__bF_buf5) );
BUFX4 BUFX4_788 ( .gnd(gnd), .vdd(vdd), .A(_4038_), .Y(_4038__bF_buf4) );
BUFX4 BUFX4_789 ( .gnd(gnd), .vdd(vdd), .A(_4038_), .Y(_4038__bF_buf3) );
BUFX4 BUFX4_790 ( .gnd(gnd), .vdd(vdd), .A(_4038_), .Y(_4038__bF_buf2) );
BUFX4 BUFX4_791 ( .gnd(gnd), .vdd(vdd), .A(_4038_), .Y(_4038__bF_buf1) );
BUFX4 BUFX4_792 ( .gnd(gnd), .vdd(vdd), .A(_4038_), .Y(_4038__bF_buf0) );
BUFX4 BUFX4_793 ( .gnd(gnd), .vdd(vdd), .A(_1031_), .Y(_1031__bF_buf3) );
BUFX4 BUFX4_794 ( .gnd(gnd), .vdd(vdd), .A(_1031_), .Y(_1031__bF_buf2) );
BUFX4 BUFX4_795 ( .gnd(gnd), .vdd(vdd), .A(_1031_), .Y(_1031__bF_buf1) );
BUFX4 BUFX4_796 ( .gnd(gnd), .vdd(vdd), .A(_1031_), .Y(_1031__bF_buf0) );
BUFX4 BUFX4_797 ( .gnd(gnd), .vdd(vdd), .A(_1507_), .Y(_1507__bF_buf7) );
BUFX4 BUFX4_798 ( .gnd(gnd), .vdd(vdd), .A(_1507_), .Y(_1507__bF_buf6) );
BUFX4 BUFX4_799 ( .gnd(gnd), .vdd(vdd), .A(_1507_), .Y(_1507__bF_buf5) );
BUFX4 BUFX4_800 ( .gnd(gnd), .vdd(vdd), .A(_1507_), .Y(_1507__bF_buf4) );
BUFX4 BUFX4_801 ( .gnd(gnd), .vdd(vdd), .A(_1507_), .Y(_1507__bF_buf3) );
BUFX4 BUFX4_802 ( .gnd(gnd), .vdd(vdd), .A(_1507_), .Y(_1507__bF_buf2) );
BUFX4 BUFX4_803 ( .gnd(gnd), .vdd(vdd), .A(_1507_), .Y(_1507__bF_buf1) );
BUFX4 BUFX4_804 ( .gnd(gnd), .vdd(vdd), .A(_1507_), .Y(_1507__bF_buf0) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf7), .B(_1104__bF_buf14), .C(regs_24__4_), .Y(_1279_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf4), .B(_1009__bF_buf3), .C(_1279_), .Y(_538_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf6), .B(_1104__bF_buf13), .C(regs_24__5_), .Y(_1280_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf3), .B(_1011__bF_buf3), .C(_1280_), .Y(_539_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf5), .B(_1104__bF_buf12), .C(regs_24__6_), .Y(_1281_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf2), .B(_1013__bF_buf3), .C(_1281_), .Y(_540_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf4), .B(_1104__bF_buf11), .C(regs_24__7_), .Y(_1282_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf1), .B(_1015__bF_buf3), .C(_1282_), .Y(_541_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf3), .B(_1104__bF_buf10), .C(regs_24__8_), .Y(_1283_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf0), .B(_1017__bF_buf3), .C(_1283_), .Y(_542_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf2), .B(_1104__bF_buf9), .C(regs_24__9_), .Y(_1284_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf4), .B(_1019__bF_buf3), .C(_1284_), .Y(_543_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf1), .B(_1104__bF_buf8), .C(regs_24__10_), .Y(_1285_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf3), .B(_1021__bF_buf3), .C(_1285_), .Y(_513_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf0), .B(_1104__bF_buf7), .C(regs_24__11_), .Y(_1286_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf2), .B(_1023__bF_buf3), .C(_1286_), .Y(_514_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf7), .B(_1104__bF_buf6), .C(regs_24__12_), .Y(_1287_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf1), .B(_1025__bF_buf3), .C(_1287_), .Y(_515_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf6), .B(_1104__bF_buf5), .C(regs_24__13_), .Y(_1288_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf0), .B(_1027__bF_buf3), .C(_1288_), .Y(_516_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf5), .B(_1104__bF_buf4), .C(regs_24__14_), .Y(_1289_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf4), .B(_1029__bF_buf3), .C(_1289_), .Y(_517_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf4), .B(_1104__bF_buf3), .C(regs_24__15_), .Y(_1290_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf3), .B(_1031__bF_buf3), .C(_1290_), .Y(_518_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf3), .B(_1104__bF_buf2), .C(regs_24__16_), .Y(_1291_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf2), .B(_1033__bF_buf3), .C(_1291_), .Y(_519_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf2), .B(_1104__bF_buf1), .C(regs_24__17_), .Y(_1292_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf1), .B(_1035__bF_buf3), .C(_1292_), .Y(_520_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf1), .B(_1104__bF_buf0), .C(regs_24__18_), .Y(_1293_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf0), .B(_1037__bF_buf3), .C(_1293_), .Y(_521_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf0), .B(_1104__bF_buf14), .C(regs_24__19_), .Y(_1294_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf4), .B(_1039__bF_buf3), .C(_1294_), .Y(_522_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf7), .B(_1104__bF_buf13), .C(regs_24__20_), .Y(_1295_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf3), .B(_1041__bF_buf3), .C(_1295_), .Y(_524_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf6), .B(_1104__bF_buf12), .C(regs_24__21_), .Y(_1296_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf2), .B(_1043__bF_buf3), .C(_1296_), .Y(_525_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf5), .B(_1104__bF_buf11), .C(regs_24__22_), .Y(_1297_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf1), .B(_1045__bF_buf3), .C(_1297_), .Y(_526_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf4), .B(_1104__bF_buf10), .C(regs_24__23_), .Y(_1298_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf0), .B(_1047__bF_buf3), .C(_1298_), .Y(_527_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf3), .B(_1104__bF_buf9), .C(regs_24__24_), .Y(_1299_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf4), .B(_1049__bF_buf3), .C(_1299_), .Y(_528_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf2), .B(_1104__bF_buf8), .C(regs_24__25_), .Y(_1300_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf3), .B(_1051__bF_buf3), .C(_1300_), .Y(_529_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf1), .B(_1104__bF_buf7), .C(regs_24__26_), .Y(_1301_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf2), .B(_1053__bF_buf3), .C(_1301_), .Y(_530_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf0), .B(_1104__bF_buf6), .C(regs_24__27_), .Y(_1302_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf1), .B(_1055__bF_buf3), .C(_1302_), .Y(_531_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf7), .B(_1104__bF_buf5), .C(regs_24__28_), .Y(_1303_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf0), .B(_1057__bF_buf3), .C(_1303_), .Y(_532_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf6), .B(_1104__bF_buf4), .C(regs_24__29_), .Y(_1304_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf4), .B(_1059__bF_buf3), .C(_1304_), .Y(_533_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf5), .B(_1104__bF_buf3), .C(regs_24__30_), .Y(_1305_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf3), .B(_1061__bF_buf3), .C(_1305_), .Y(_535_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf4), .B(_1104__bF_buf2), .C(regs_24__31_), .Y(_1306_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf2), .B(_1063__bF_buf3), .C(_1306_), .Y(_536_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(regs_23__0_), .Y(_1307_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(waddr[3]), .B(_993_), .Y(_1308_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_1308_), .B(waddr[2]), .Y(_1309_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_1142__bF_buf5), .B(_1309__bF_buf5), .Y(_1310_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(wdata[0]), .B(_1310__bF_buf7), .Y(_1311_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1307_), .B(_1310__bF_buf6), .C(_1311_), .Y(_480_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(regs_23__1_), .Y(_1312_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(wdata[1]), .B(_1310__bF_buf5), .Y(_1313_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1312_), .B(_1310__bF_buf4), .C(_1313_), .Y(_491_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(regs_23__2_), .Y(_1314_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(wdata[2]), .B(_1310__bF_buf3), .Y(_1315_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1314_), .B(_1310__bF_buf2), .C(_1315_), .Y(_502_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(regs_23__3_), .Y(_1316_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(wdata[3]), .B(_1310__bF_buf1), .Y(_1317_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1316_), .B(_1310__bF_buf0), .C(_1317_), .Y(_505_) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(regs_23__4_), .Y(_1318_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(wdata[4]), .B(_1310__bF_buf7), .Y(_1319_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1318_), .B(_1310__bF_buf6), .C(_1319_), .Y(_506_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(regs_23__5_), .Y(_1320_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(wdata[5]), .B(_1310__bF_buf5), .Y(_1321_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1320_), .B(_1310__bF_buf4), .C(_1321_), .Y(_507_) );
INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(regs_23__6_), .Y(_1322_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(wdata[6]), .B(_1310__bF_buf3), .Y(_1323_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1322_), .B(_1310__bF_buf2), .C(_1323_), .Y(_508_) );
INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(regs_23__7_), .Y(_1324_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(wdata[7]), .B(_1310__bF_buf1), .Y(_1325_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1324_), .B(_1310__bF_buf0), .C(_1325_), .Y(_509_) );
INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(regs_23__8_), .Y(_1326_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(wdata[8]), .B(_1310__bF_buf7), .Y(_1327_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_1326_), .B(_1310__bF_buf6), .C(_1327_), .Y(_510_) );
INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(regs_23__9_), .Y(_1328_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(wdata[9]), .B(_1310__bF_buf5), .Y(_1329_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_1328_), .B(_1310__bF_buf4), .C(_1329_), .Y(_511_) );
INVX2 INVX2_11 ( .gnd(gnd), .vdd(vdd), .A(regs_23__10_), .Y(_1330_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(wdata[10]), .B(_1310__bF_buf3), .Y(_1331_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_1330_), .B(_1310__bF_buf2), .C(_1331_), .Y(_481_) );
INVX2 INVX2_12 ( .gnd(gnd), .vdd(vdd), .A(regs_23__11_), .Y(_1332_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(wdata[11]), .B(_1310__bF_buf1), .Y(_1333_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1332_), .B(_1310__bF_buf0), .C(_1333_), .Y(_482_) );
INVX2 INVX2_13 ( .gnd(gnd), .vdd(vdd), .A(regs_23__12_), .Y(_1334_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(wdata[12]), .B(_1310__bF_buf7), .Y(_1335_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_1334_), .B(_1310__bF_buf6), .C(_1335_), .Y(_483_) );
INVX2 INVX2_14 ( .gnd(gnd), .vdd(vdd), .A(regs_23__13_), .Y(_1336_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(wdata[13]), .B(_1310__bF_buf5), .Y(_1337_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_1336_), .B(_1310__bF_buf4), .C(_1337_), .Y(_484_) );
INVX2 INVX2_15 ( .gnd(gnd), .vdd(vdd), .A(regs_23__14_), .Y(_1338_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(wdata[14]), .B(_1310__bF_buf3), .Y(_1339_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1338_), .B(_1310__bF_buf2), .C(_1339_), .Y(_485_) );
INVX2 INVX2_16 ( .gnd(gnd), .vdd(vdd), .A(regs_23__15_), .Y(_1340_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(wdata[15]), .B(_1310__bF_buf1), .Y(_1341_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1340_), .B(_1310__bF_buf0), .C(_1341_), .Y(_486_) );
INVX2 INVX2_17 ( .gnd(gnd), .vdd(vdd), .A(regs_23__16_), .Y(_1342_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(wdata[16]), .B(_1310__bF_buf7), .Y(_1343_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1342_), .B(_1310__bF_buf6), .C(_1343_), .Y(_487_) );
INVX2 INVX2_18 ( .gnd(gnd), .vdd(vdd), .A(regs_23__17_), .Y(_1344_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(wdata[17]), .B(_1310__bF_buf5), .Y(_1345_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_1344_), .B(_1310__bF_buf4), .C(_1345_), .Y(_488_) );
INVX2 INVX2_19 ( .gnd(gnd), .vdd(vdd), .A(regs_23__18_), .Y(_1346_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(wdata[18]), .B(_1310__bF_buf3), .Y(_1347_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_1346_), .B(_1310__bF_buf2), .C(_1347_), .Y(_489_) );
INVX2 INVX2_20 ( .gnd(gnd), .vdd(vdd), .A(regs_23__19_), .Y(_1348_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(wdata[19]), .B(_1310__bF_buf1), .Y(_1349_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_1348_), .B(_1310__bF_buf0), .C(_1349_), .Y(_490_) );
INVX2 INVX2_21 ( .gnd(gnd), .vdd(vdd), .A(regs_23__20_), .Y(_1350_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(wdata[20]), .B(_1310__bF_buf7), .Y(_1351_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_1350_), .B(_1310__bF_buf6), .C(_1351_), .Y(_492_) );
INVX2 INVX2_22 ( .gnd(gnd), .vdd(vdd), .A(regs_23__21_), .Y(_1352_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(wdata[21]), .B(_1310__bF_buf5), .Y(_1353_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1352_), .B(_1310__bF_buf4), .C(_1353_), .Y(_493_) );
INVX2 INVX2_23 ( .gnd(gnd), .vdd(vdd), .A(regs_23__22_), .Y(_1354_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(wdata[22]), .B(_1310__bF_buf3), .Y(_1355_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_1354_), .B(_1310__bF_buf2), .C(_1355_), .Y(_494_) );
INVX2 INVX2_24 ( .gnd(gnd), .vdd(vdd), .A(regs_23__23_), .Y(_1356_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(wdata[23]), .B(_1310__bF_buf1), .Y(_1357_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_1356_), .B(_1310__bF_buf0), .C(_1357_), .Y(_495_) );
INVX2 INVX2_25 ( .gnd(gnd), .vdd(vdd), .A(regs_23__24_), .Y(_1358_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(wdata[24]), .B(_1310__bF_buf7), .Y(_1359_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1358_), .B(_1310__bF_buf6), .C(_1359_), .Y(_496_) );
INVX2 INVX2_26 ( .gnd(gnd), .vdd(vdd), .A(regs_23__25_), .Y(_1360_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(wdata[25]), .B(_1310__bF_buf5), .Y(_1361_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1360_), .B(_1310__bF_buf4), .C(_1361_), .Y(_497_) );
INVX2 INVX2_27 ( .gnd(gnd), .vdd(vdd), .A(regs_23__26_), .Y(_1362_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(wdata[26]), .B(_1310__bF_buf3), .Y(_1363_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1362_), .B(_1310__bF_buf2), .C(_1363_), .Y(_498_) );
INVX2 INVX2_28 ( .gnd(gnd), .vdd(vdd), .A(regs_23__27_), .Y(_1364_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(wdata[27]), .B(_1310__bF_buf1), .Y(_1365_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_1364_), .B(_1310__bF_buf0), .C(_1365_), .Y(_499_) );
INVX2 INVX2_29 ( .gnd(gnd), .vdd(vdd), .A(regs_23__28_), .Y(_1366_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(wdata[28]), .B(_1310__bF_buf7), .Y(_1367_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1366_), .B(_1310__bF_buf6), .C(_1367_), .Y(_500_) );
INVX2 INVX2_30 ( .gnd(gnd), .vdd(vdd), .A(regs_23__29_), .Y(_1368_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(wdata[29]), .B(_1310__bF_buf5), .Y(_1369_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1368_), .B(_1310__bF_buf4), .C(_1369_), .Y(_501_) );
INVX2 INVX2_31 ( .gnd(gnd), .vdd(vdd), .A(regs_23__30_), .Y(_1370_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(wdata[30]), .B(_1310__bF_buf3), .Y(_1371_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1370_), .B(_1310__bF_buf2), .C(_1371_), .Y(_503_) );
INVX2 INVX2_32 ( .gnd(gnd), .vdd(vdd), .A(regs_23__31_), .Y(_1372_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(wdata[31]), .B(_1310__bF_buf1), .Y(_1373_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1372_), .B(_1310__bF_buf0), .C(_1373_), .Y(_504_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf9), .B(_1309__bF_buf4), .Y(_1374_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(regs_22__0_), .B(_1374__bF_buf7), .Y(_1375_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_992__bF_buf3), .B(_1374__bF_buf6), .C(_1375_), .Y(_448_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(regs_22__1_), .B(_1374__bF_buf5), .Y(_1376_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_1003__bF_buf3), .B(_1374__bF_buf4), .C(_1376_), .Y(_459_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(regs_22__2_), .B(_1374__bF_buf3), .Y(_1377_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf3), .B(_1374__bF_buf2), .C(_1377_), .Y(_470_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(regs_22__3_), .B(_1374__bF_buf1), .Y(_1378_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_1007__bF_buf3), .B(_1374__bF_buf0), .C(_1378_), .Y(_473_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(regs_22__4_), .B(_1374__bF_buf7), .Y(_1379_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_1009__bF_buf2), .B(_1374__bF_buf6), .C(_1379_), .Y(_474_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(regs_22__5_), .B(_1374__bF_buf5), .Y(_1380_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_1011__bF_buf2), .B(_1374__bF_buf4), .C(_1380_), .Y(_475_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(regs_22__6_), .B(_1374__bF_buf3), .Y(_1381_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1013__bF_buf2), .B(_1374__bF_buf2), .C(_1381_), .Y(_476_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(regs_22__7_), .B(_1374__bF_buf1), .Y(_1382_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_1015__bF_buf2), .B(_1374__bF_buf0), .C(_1382_), .Y(_477_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(regs_22__8_), .B(_1374__bF_buf7), .Y(_1383_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf2), .B(_1374__bF_buf6), .C(_1383_), .Y(_478_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(regs_22__9_), .B(_1374__bF_buf5), .Y(_1384_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_1019__bF_buf2), .B(_1374__bF_buf4), .C(_1384_), .Y(_479_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(regs_22__10_), .B(_1374__bF_buf3), .Y(_1385_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1021__bF_buf2), .B(_1374__bF_buf2), .C(_1385_), .Y(_449_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(regs_22__11_), .B(_1374__bF_buf1), .Y(_1386_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1023__bF_buf2), .B(_1374__bF_buf0), .C(_1386_), .Y(_450_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(regs_22__12_), .B(_1374__bF_buf7), .Y(_1387_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1025__bF_buf2), .B(_1374__bF_buf6), .C(_1387_), .Y(_451_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(regs_22__13_), .B(_1374__bF_buf5), .Y(_1388_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_1027__bF_buf2), .B(_1374__bF_buf4), .C(_1388_), .Y(_452_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(regs_22__14_), .B(_1374__bF_buf3), .Y(_1389_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1029__bF_buf2), .B(_1374__bF_buf2), .C(_1389_), .Y(_453_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(regs_22__15_), .B(_1374__bF_buf1), .Y(_1390_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf2), .B(_1374__bF_buf0), .C(_1390_), .Y(_454_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(regs_22__16_), .B(_1374__bF_buf7), .Y(_1391_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1033__bF_buf2), .B(_1374__bF_buf6), .C(_1391_), .Y(_455_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(regs_22__17_), .B(_1374__bF_buf5), .Y(_1392_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1035__bF_buf2), .B(_1374__bF_buf4), .C(_1392_), .Y(_456_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(regs_22__18_), .B(_1374__bF_buf3), .Y(_1393_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1037__bF_buf2), .B(_1374__bF_buf2), .C(_1393_), .Y(_457_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(regs_22__19_), .B(_1374__bF_buf1), .Y(_1394_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1039__bF_buf2), .B(_1374__bF_buf0), .C(_1394_), .Y(_458_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(regs_22__20_), .B(_1374__bF_buf7), .Y(_1395_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_1041__bF_buf2), .B(_1374__bF_buf6), .C(_1395_), .Y(_460_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(regs_22__21_), .B(_1374__bF_buf5), .Y(_1396_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_1043__bF_buf2), .B(_1374__bF_buf4), .C(_1396_), .Y(_461_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(regs_22__22_), .B(_1374__bF_buf3), .Y(_1397_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_1045__bF_buf2), .B(_1374__bF_buf2), .C(_1397_), .Y(_462_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(regs_22__23_), .B(_1374__bF_buf1), .Y(_1398_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_1047__bF_buf2), .B(_1374__bF_buf0), .C(_1398_), .Y(_463_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(regs_22__24_), .B(_1374__bF_buf7), .Y(_1399_) );
AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1049__bF_buf2), .B(_1374__bF_buf6), .C(_1399_), .Y(_464_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(regs_22__25_), .B(_1374__bF_buf5), .Y(_1400_) );
AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_1051__bF_buf2), .B(_1374__bF_buf4), .C(_1400_), .Y(_465_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(regs_22__26_), .B(_1374__bF_buf3), .Y(_1401_) );
AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1053__bF_buf2), .B(_1374__bF_buf2), .C(_1401_), .Y(_466_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(regs_22__27_), .B(_1374__bF_buf1), .Y(_1402_) );
AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_1055__bF_buf2), .B(_1374__bF_buf0), .C(_1402_), .Y(_467_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(regs_22__28_), .B(_1374__bF_buf7), .Y(_1403_) );
AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_1057__bF_buf2), .B(_1374__bF_buf6), .C(_1403_), .Y(_468_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(regs_22__29_), .B(_1374__bF_buf5), .Y(_1404_) );
AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_1059__bF_buf2), .B(_1374__bF_buf4), .C(_1404_), .Y(_469_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(regs_22__30_), .B(_1374__bF_buf3), .Y(_1405_) );
AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1061__bF_buf2), .B(_1374__bF_buf2), .C(_1405_), .Y(_471_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(regs_22__31_), .B(_1374__bF_buf1), .Y(_1406_) );
AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1063__bF_buf2), .B(_1374__bF_buf0), .C(_1406_), .Y(_472_) );
INVX2 INVX2_33 ( .gnd(gnd), .vdd(vdd), .A(regs_21__0_), .Y(_1407_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf3), .B(_1070__bF_buf10), .Y(_1408_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(wdata[0]), .B(_1408__bF_buf7), .Y(_1409_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1407_), .B(_1408__bF_buf6), .C(_1409_), .Y(_416_) );
INVX2 INVX2_34 ( .gnd(gnd), .vdd(vdd), .A(regs_21__1_), .Y(_1410_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(wdata[1]), .B(_1408__bF_buf5), .Y(_1411_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1410_), .B(_1408__bF_buf4), .C(_1411_), .Y(_427_) );
INVX2 INVX2_35 ( .gnd(gnd), .vdd(vdd), .A(regs_21__2_), .Y(_1412_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(wdata[2]), .B(_1408__bF_buf3), .Y(_1413_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1412_), .B(_1408__bF_buf2), .C(_1413_), .Y(_438_) );
INVX2 INVX2_36 ( .gnd(gnd), .vdd(vdd), .A(regs_21__3_), .Y(_1414_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(wdata[3]), .B(_1408__bF_buf1), .Y(_1415_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1414_), .B(_1408__bF_buf0), .C(_1415_), .Y(_441_) );
INVX2 INVX2_37 ( .gnd(gnd), .vdd(vdd), .A(regs_21__4_), .Y(_1416_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(wdata[4]), .B(_1408__bF_buf7), .Y(_1417_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_1416_), .B(_1408__bF_buf6), .C(_1417_), .Y(_442_) );
INVX2 INVX2_38 ( .gnd(gnd), .vdd(vdd), .A(regs_21__5_), .Y(_1418_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(wdata[5]), .B(_1408__bF_buf5), .Y(_1419_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1418_), .B(_1408__bF_buf4), .C(_1419_), .Y(_443_) );
INVX2 INVX2_39 ( .gnd(gnd), .vdd(vdd), .A(regs_21__6_), .Y(_1420_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(wdata[6]), .B(_1408__bF_buf3), .Y(_1421_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(_1408__bF_buf2), .C(_1421_), .Y(_444_) );
INVX2 INVX2_40 ( .gnd(gnd), .vdd(vdd), .A(regs_21__7_), .Y(_1422_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(wdata[7]), .B(_1408__bF_buf1), .Y(_1423_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1422_), .B(_1408__bF_buf0), .C(_1423_), .Y(_445_) );
INVX2 INVX2_41 ( .gnd(gnd), .vdd(vdd), .A(regs_21__8_), .Y(_1424_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(wdata[8]), .B(_1408__bF_buf7), .Y(_1425_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1424_), .B(_1408__bF_buf6), .C(_1425_), .Y(_446_) );
INVX2 INVX2_42 ( .gnd(gnd), .vdd(vdd), .A(regs_21__9_), .Y(_1426_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(wdata[9]), .B(_1408__bF_buf5), .Y(_1427_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1426_), .B(_1408__bF_buf4), .C(_1427_), .Y(_447_) );
INVX2 INVX2_43 ( .gnd(gnd), .vdd(vdd), .A(regs_21__10_), .Y(_1428_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(wdata[10]), .B(_1408__bF_buf3), .Y(_1429_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1428_), .B(_1408__bF_buf2), .C(_1429_), .Y(_417_) );
INVX2 INVX2_44 ( .gnd(gnd), .vdd(vdd), .A(regs_21__11_), .Y(_1430_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(wdata[11]), .B(_1408__bF_buf1), .Y(_1431_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1430_), .B(_1408__bF_buf0), .C(_1431_), .Y(_418_) );
INVX2 INVX2_45 ( .gnd(gnd), .vdd(vdd), .A(regs_21__12_), .Y(_1432_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(wdata[12]), .B(_1408__bF_buf7), .Y(_1433_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1432_), .B(_1408__bF_buf6), .C(_1433_), .Y(_419_) );
INVX2 INVX2_46 ( .gnd(gnd), .vdd(vdd), .A(regs_21__13_), .Y(_1434_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(wdata[13]), .B(_1408__bF_buf5), .Y(_1435_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1434_), .B(_1408__bF_buf4), .C(_1435_), .Y(_420_) );
INVX2 INVX2_47 ( .gnd(gnd), .vdd(vdd), .A(regs_21__14_), .Y(_1436_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(wdata[14]), .B(_1408__bF_buf3), .Y(_1437_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1436_), .B(_1408__bF_buf2), .C(_1437_), .Y(_421_) );
INVX2 INVX2_48 ( .gnd(gnd), .vdd(vdd), .A(regs_21__15_), .Y(_1438_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(wdata[15]), .B(_1408__bF_buf1), .Y(_1439_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1438_), .B(_1408__bF_buf0), .C(_1439_), .Y(_422_) );
INVX2 INVX2_49 ( .gnd(gnd), .vdd(vdd), .A(regs_21__16_), .Y(_1440_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(wdata[16]), .B(_1408__bF_buf7), .Y(_1441_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1440_), .B(_1408__bF_buf6), .C(_1441_), .Y(_423_) );
INVX2 INVX2_50 ( .gnd(gnd), .vdd(vdd), .A(regs_21__17_), .Y(_1442_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(wdata[17]), .B(_1408__bF_buf5), .Y(_1443_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1442_), .B(_1408__bF_buf4), .C(_1443_), .Y(_424_) );
INVX2 INVX2_51 ( .gnd(gnd), .vdd(vdd), .A(regs_21__18_), .Y(_1444_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(wdata[18]), .B(_1408__bF_buf3), .Y(_1445_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1444_), .B(_1408__bF_buf2), .C(_1445_), .Y(_425_) );
INVX2 INVX2_52 ( .gnd(gnd), .vdd(vdd), .A(regs_21__19_), .Y(_1446_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(wdata[19]), .B(_1408__bF_buf1), .Y(_1447_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_1446_), .B(_1408__bF_buf0), .C(_1447_), .Y(_426_) );
INVX2 INVX2_53 ( .gnd(gnd), .vdd(vdd), .A(regs_21__20_), .Y(_1448_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(wdata[20]), .B(_1408__bF_buf7), .Y(_1449_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1448_), .B(_1408__bF_buf6), .C(_1449_), .Y(_428_) );
INVX2 INVX2_54 ( .gnd(gnd), .vdd(vdd), .A(regs_21__21_), .Y(_1450_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(wdata[21]), .B(_1408__bF_buf5), .Y(_1451_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1450_), .B(_1408__bF_buf4), .C(_1451_), .Y(_429_) );
INVX2 INVX2_55 ( .gnd(gnd), .vdd(vdd), .A(regs_21__22_), .Y(_1452_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(wdata[22]), .B(_1408__bF_buf3), .Y(_1453_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1452_), .B(_1408__bF_buf2), .C(_1453_), .Y(_430_) );
INVX2 INVX2_56 ( .gnd(gnd), .vdd(vdd), .A(regs_21__23_), .Y(_1454_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(wdata[23]), .B(_1408__bF_buf1), .Y(_1455_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1454_), .B(_1408__bF_buf0), .C(_1455_), .Y(_431_) );
INVX2 INVX2_57 ( .gnd(gnd), .vdd(vdd), .A(regs_21__24_), .Y(_1456_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(wdata[24]), .B(_1408__bF_buf7), .Y(_1457_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1456_), .B(_1408__bF_buf6), .C(_1457_), .Y(_432_) );
INVX2 INVX2_58 ( .gnd(gnd), .vdd(vdd), .A(regs_21__25_), .Y(_1458_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(wdata[25]), .B(_1408__bF_buf5), .Y(_1459_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1458_), .B(_1408__bF_buf4), .C(_1459_), .Y(_433_) );
INVX2 INVX2_59 ( .gnd(gnd), .vdd(vdd), .A(regs_21__26_), .Y(_1460_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(wdata[26]), .B(_1408__bF_buf3), .Y(_1461_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_1460_), .B(_1408__bF_buf2), .C(_1461_), .Y(_434_) );
INVX2 INVX2_60 ( .gnd(gnd), .vdd(vdd), .A(regs_21__27_), .Y(_1462_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(wdata[27]), .B(_1408__bF_buf1), .Y(_1463_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1462_), .B(_1408__bF_buf0), .C(_1463_), .Y(_435_) );
INVX2 INVX2_61 ( .gnd(gnd), .vdd(vdd), .A(regs_21__28_), .Y(_1464_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(wdata[28]), .B(_1408__bF_buf7), .Y(_1465_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(_1408__bF_buf6), .C(_1465_), .Y(_436_) );
INVX2 INVX2_62 ( .gnd(gnd), .vdd(vdd), .A(regs_21__29_), .Y(_1466_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(wdata[29]), .B(_1408__bF_buf5), .Y(_1467_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1466_), .B(_1408__bF_buf4), .C(_1467_), .Y(_437_) );
INVX2 INVX2_63 ( .gnd(gnd), .vdd(vdd), .A(regs_21__30_), .Y(_1468_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(wdata[30]), .B(_1408__bF_buf3), .Y(_1469_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1468_), .B(_1408__bF_buf2), .C(_1469_), .Y(_439_) );
INVX2 INVX2_64 ( .gnd(gnd), .vdd(vdd), .A(regs_21__31_), .Y(_1470_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(wdata[31]), .B(_1408__bF_buf1), .Y(_1471_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1470_), .B(_1408__bF_buf0), .C(_1471_), .Y(_440_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf2), .B(_1104__bF_buf1), .Y(_1472_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf1), .B(_1104__bF_buf0), .C(regs_20__0_), .Y(_1473_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf4), .B(_992__bF_buf2), .C(_1473_), .Y(_384_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf0), .B(_1104__bF_buf14), .C(regs_20__1_), .Y(_1474_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf3), .B(_1003__bF_buf2), .C(_1474_), .Y(_395_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf5), .B(_1104__bF_buf13), .C(regs_20__2_), .Y(_1475_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf2), .B(_1005__bF_buf2), .C(_1475_), .Y(_406_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf4), .B(_1104__bF_buf12), .C(regs_20__3_), .Y(_1476_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf1), .B(_1007__bF_buf2), .C(_1476_), .Y(_409_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf3), .B(_1104__bF_buf11), .C(regs_20__4_), .Y(_1477_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf0), .B(_1009__bF_buf1), .C(_1477_), .Y(_410_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf2), .B(_1104__bF_buf10), .C(regs_20__5_), .Y(_1478_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf4), .B(_1011__bF_buf1), .C(_1478_), .Y(_411_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf1), .B(_1104__bF_buf9), .C(regs_20__6_), .Y(_1479_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf3), .B(_1013__bF_buf1), .C(_1479_), .Y(_412_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf0), .B(_1104__bF_buf8), .C(regs_20__7_), .Y(_1480_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf2), .B(_1015__bF_buf1), .C(_1480_), .Y(_413_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf5), .B(_1104__bF_buf7), .C(regs_20__8_), .Y(_1481_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf1), .B(_1017__bF_buf1), .C(_1481_), .Y(_414_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf4), .B(_1104__bF_buf6), .C(regs_20__9_), .Y(_1482_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf0), .B(_1019__bF_buf1), .C(_1482_), .Y(_415_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf3), .B(_1104__bF_buf5), .C(regs_20__10_), .Y(_1483_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf4), .B(_1021__bF_buf1), .C(_1483_), .Y(_385_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf2), .B(_1104__bF_buf4), .C(regs_20__11_), .Y(_1484_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf3), .B(_1023__bF_buf1), .C(_1484_), .Y(_386_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf1), .B(_1104__bF_buf3), .C(regs_20__12_), .Y(_1485_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf2), .B(_1025__bF_buf1), .C(_1485_), .Y(_387_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf0), .B(_1104__bF_buf2), .C(regs_20__13_), .Y(_1486_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf1), .B(_1027__bF_buf1), .C(_1486_), .Y(_388_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf5), .B(_1104__bF_buf1), .C(regs_20__14_), .Y(_1487_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf0), .B(_1029__bF_buf1), .C(_1487_), .Y(_389_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf4), .B(_1104__bF_buf0), .C(regs_20__15_), .Y(_1488_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf4), .B(_1031__bF_buf1), .C(_1488_), .Y(_390_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf3), .B(_1104__bF_buf14), .C(regs_20__16_), .Y(_1489_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf3), .B(_1033__bF_buf1), .C(_1489_), .Y(_391_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf2), .B(_1104__bF_buf13), .C(regs_20__17_), .Y(_1490_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf2), .B(_1035__bF_buf1), .C(_1490_), .Y(_392_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf1), .B(_1104__bF_buf12), .C(regs_20__18_), .Y(_1491_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf1), .B(_1037__bF_buf1), .C(_1491_), .Y(_393_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf0), .B(_1104__bF_buf11), .C(regs_20__19_), .Y(_1492_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf0), .B(_1039__bF_buf1), .C(_1492_), .Y(_394_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf5), .B(_1104__bF_buf10), .C(regs_20__20_), .Y(_1493_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf4), .B(_1041__bF_buf1), .C(_1493_), .Y(_396_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf4), .B(_1104__bF_buf9), .C(regs_20__21_), .Y(_1494_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf3), .B(_1043__bF_buf1), .C(_1494_), .Y(_397_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf3), .B(_1104__bF_buf8), .C(regs_20__22_), .Y(_1495_) );
OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf2), .B(_1045__bF_buf1), .C(_1495_), .Y(_398_) );
OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf2), .B(_1104__bF_buf7), .C(regs_20__23_), .Y(_1496_) );
OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf1), .B(_1047__bF_buf1), .C(_1496_), .Y(_399_) );
OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf1), .B(_1104__bF_buf6), .C(regs_20__24_), .Y(_1497_) );
OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf0), .B(_1049__bF_buf1), .C(_1497_), .Y(_400_) );
OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf0), .B(_1104__bF_buf5), .C(regs_20__25_), .Y(_1498_) );
OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf4), .B(_1051__bF_buf1), .C(_1498_), .Y(_401_) );
OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf5), .B(_1104__bF_buf4), .C(regs_20__26_), .Y(_1499_) );
OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf3), .B(_1053__bF_buf1), .C(_1499_), .Y(_402_) );
OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf4), .B(_1104__bF_buf3), .C(regs_20__27_), .Y(_1500_) );
OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf2), .B(_1055__bF_buf1), .C(_1500_), .Y(_403_) );
OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf3), .B(_1104__bF_buf2), .C(regs_20__28_), .Y(_1501_) );
OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf1), .B(_1057__bF_buf1), .C(_1501_), .Y(_404_) );
OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf2), .B(_1104__bF_buf1), .C(regs_20__29_), .Y(_1502_) );
OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf0), .B(_1059__bF_buf1), .C(_1502_), .Y(_405_) );
OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf1), .B(_1104__bF_buf0), .C(regs_20__30_), .Y(_1503_) );
OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf4), .B(_1061__bF_buf1), .C(_1503_), .Y(_407_) );
OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1309__bF_buf0), .B(_1104__bF_buf14), .C(regs_20__31_), .Y(_1504_) );
OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_1472__bF_buf3), .B(_1063__bF_buf1), .C(_1504_), .Y(_408_) );
INVX2 INVX2_65 ( .gnd(gnd), .vdd(vdd), .A(regs_19__0_), .Y(_1505_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_1308_), .B(_1139_), .Y(_1506_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1142__bF_buf4), .B(_1506__bF_buf5), .Y(_1507_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(wdata[0]), .B(_1507__bF_buf7), .Y(_1508_) );
OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1505_), .B(_1507__bF_buf6), .C(_1508_), .Y(_320_) );
INVX2 INVX2_66 ( .gnd(gnd), .vdd(vdd), .A(regs_19__1_), .Y(_1509_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(wdata[1]), .B(_1507__bF_buf5), .Y(_1510_) );
OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_1509_), .B(_1507__bF_buf4), .C(_1510_), .Y(_331_) );
INVX2 INVX2_67 ( .gnd(gnd), .vdd(vdd), .A(regs_19__2_), .Y(_1511_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(wdata[2]), .B(_1507__bF_buf3), .Y(_1512_) );
OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1511_), .B(_1507__bF_buf2), .C(_1512_), .Y(_342_) );
INVX2 INVX2_68 ( .gnd(gnd), .vdd(vdd), .A(regs_19__3_), .Y(_1513_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(wdata[3]), .B(_1507__bF_buf1), .Y(_1514_) );
OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1513_), .B(_1507__bF_buf0), .C(_1514_), .Y(_345_) );
INVX2 INVX2_69 ( .gnd(gnd), .vdd(vdd), .A(regs_19__4_), .Y(_1515_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(wdata[4]), .B(_1507__bF_buf7), .Y(_1516_) );
OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1515_), .B(_1507__bF_buf6), .C(_1516_), .Y(_346_) );
INVX2 INVX2_70 ( .gnd(gnd), .vdd(vdd), .A(regs_19__5_), .Y(_1517_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(wdata[5]), .B(_1507__bF_buf5), .Y(_1518_) );
OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1517_), .B(_1507__bF_buf4), .C(_1518_), .Y(_347_) );
INVX2 INVX2_71 ( .gnd(gnd), .vdd(vdd), .A(regs_19__6_), .Y(_1519_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(wdata[6]), .B(_1507__bF_buf3), .Y(_1520_) );
OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1519_), .B(_1507__bF_buf2), .C(_1520_), .Y(_348_) );
INVX2 INVX2_72 ( .gnd(gnd), .vdd(vdd), .A(regs_19__7_), .Y(_1521_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(wdata[7]), .B(_1507__bF_buf1), .Y(_1522_) );
OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1521_), .B(_1507__bF_buf0), .C(_1522_), .Y(_349_) );
INVX2 INVX2_73 ( .gnd(gnd), .vdd(vdd), .A(regs_19__8_), .Y(_1523_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(wdata[8]), .B(_1507__bF_buf7), .Y(_1524_) );
OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1523_), .B(_1507__bF_buf6), .C(_1524_), .Y(_350_) );
INVX2 INVX2_74 ( .gnd(gnd), .vdd(vdd), .A(regs_19__9_), .Y(_1525_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(wdata[9]), .B(_1507__bF_buf5), .Y(_1526_) );
OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1525_), .B(_1507__bF_buf4), .C(_1526_), .Y(_351_) );
INVX2 INVX2_75 ( .gnd(gnd), .vdd(vdd), .A(regs_19__10_), .Y(_1527_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(wdata[10]), .B(_1507__bF_buf3), .Y(_1528_) );
OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1527_), .B(_1507__bF_buf2), .C(_1528_), .Y(_321_) );
INVX2 INVX2_76 ( .gnd(gnd), .vdd(vdd), .A(regs_19__11_), .Y(_1529_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(wdata[11]), .B(_1507__bF_buf1), .Y(_1530_) );
OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1529_), .B(_1507__bF_buf0), .C(_1530_), .Y(_322_) );
INVX2 INVX2_77 ( .gnd(gnd), .vdd(vdd), .A(regs_19__12_), .Y(_1531_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(wdata[12]), .B(_1507__bF_buf7), .Y(_1532_) );
OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1531_), .B(_1507__bF_buf6), .C(_1532_), .Y(_323_) );
INVX2 INVX2_78 ( .gnd(gnd), .vdd(vdd), .A(regs_19__13_), .Y(_1533_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(wdata[13]), .B(_1507__bF_buf5), .Y(_1534_) );
OAI21X1 OAI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1533_), .B(_1507__bF_buf4), .C(_1534_), .Y(_324_) );
INVX2 INVX2_79 ( .gnd(gnd), .vdd(vdd), .A(regs_19__14_), .Y(_1535_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(wdata[14]), .B(_1507__bF_buf3), .Y(_1536_) );
OAI21X1 OAI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1535_), .B(_1507__bF_buf2), .C(_1536_), .Y(_325_) );
INVX2 INVX2_80 ( .gnd(gnd), .vdd(vdd), .A(regs_19__15_), .Y(_1537_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(wdata[15]), .B(_1507__bF_buf1), .Y(_1538_) );
OAI21X1 OAI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1537_), .B(_1507__bF_buf0), .C(_1538_), .Y(_326_) );
INVX2 INVX2_81 ( .gnd(gnd), .vdd(vdd), .A(regs_19__16_), .Y(_1539_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(wdata[16]), .B(_1507__bF_buf7), .Y(_1540_) );
OAI21X1 OAI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1539_), .B(_1507__bF_buf6), .C(_1540_), .Y(_327_) );
INVX2 INVX2_82 ( .gnd(gnd), .vdd(vdd), .A(regs_19__17_), .Y(_1541_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(wdata[17]), .B(_1507__bF_buf5), .Y(_1542_) );
OAI21X1 OAI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1541_), .B(_1507__bF_buf4), .C(_1542_), .Y(_328_) );
INVX2 INVX2_83 ( .gnd(gnd), .vdd(vdd), .A(regs_19__18_), .Y(_1543_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(wdata[18]), .B(_1507__bF_buf3), .Y(_1544_) );
OAI21X1 OAI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1543_), .B(_1507__bF_buf2), .C(_1544_), .Y(_329_) );
INVX2 INVX2_84 ( .gnd(gnd), .vdd(vdd), .A(regs_19__19_), .Y(_1545_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(wdata[19]), .B(_1507__bF_buf1), .Y(_1546_) );
OAI21X1 OAI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_1545_), .B(_1507__bF_buf0), .C(_1546_), .Y(_330_) );
INVX2 INVX2_85 ( .gnd(gnd), .vdd(vdd), .A(regs_19__20_), .Y(_1547_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(wdata[20]), .B(_1507__bF_buf7), .Y(_1548_) );
OAI21X1 OAI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_1547_), .B(_1507__bF_buf6), .C(_1548_), .Y(_332_) );
INVX2 INVX2_86 ( .gnd(gnd), .vdd(vdd), .A(regs_19__21_), .Y(_1549_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(wdata[21]), .B(_1507__bF_buf5), .Y(_1550_) );
OAI21X1 OAI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1549_), .B(_1507__bF_buf4), .C(_1550_), .Y(_333_) );
INVX2 INVX2_87 ( .gnd(gnd), .vdd(vdd), .A(regs_19__22_), .Y(_1551_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(wdata[22]), .B(_1507__bF_buf3), .Y(_1552_) );
OAI21X1 OAI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1551_), .B(_1507__bF_buf2), .C(_1552_), .Y(_334_) );
INVX2 INVX2_88 ( .gnd(gnd), .vdd(vdd), .A(regs_19__23_), .Y(_1553_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(wdata[23]), .B(_1507__bF_buf1), .Y(_1554_) );
OAI21X1 OAI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_1553_), .B(_1507__bF_buf0), .C(_1554_), .Y(_335_) );
INVX2 INVX2_89 ( .gnd(gnd), .vdd(vdd), .A(regs_19__24_), .Y(_1555_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(wdata[24]), .B(_1507__bF_buf7), .Y(_1556_) );
OAI21X1 OAI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1555_), .B(_1507__bF_buf6), .C(_1556_), .Y(_336_) );
INVX2 INVX2_90 ( .gnd(gnd), .vdd(vdd), .A(regs_19__25_), .Y(_1557_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(wdata[25]), .B(_1507__bF_buf5), .Y(_1558_) );
OAI21X1 OAI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1557_), .B(_1507__bF_buf4), .C(_1558_), .Y(_337_) );
INVX2 INVX2_91 ( .gnd(gnd), .vdd(vdd), .A(regs_19__26_), .Y(_1559_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(wdata[26]), .B(_1507__bF_buf3), .Y(_1560_) );
OAI21X1 OAI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1559_), .B(_1507__bF_buf2), .C(_1560_), .Y(_338_) );
INVX2 INVX2_92 ( .gnd(gnd), .vdd(vdd), .A(regs_19__27_), .Y(_1561_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(wdata[27]), .B(_1507__bF_buf1), .Y(_1562_) );
OAI21X1 OAI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .B(_1507__bF_buf0), .C(_1562_), .Y(_339_) );
INVX2 INVX2_93 ( .gnd(gnd), .vdd(vdd), .A(regs_19__28_), .Y(_1563_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(wdata[28]), .B(_1507__bF_buf7), .Y(_1564_) );
OAI21X1 OAI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1563_), .B(_1507__bF_buf6), .C(_1564_), .Y(_340_) );
INVX2 INVX2_94 ( .gnd(gnd), .vdd(vdd), .A(regs_19__29_), .Y(_1565_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(wdata[29]), .B(_1507__bF_buf5), .Y(_1566_) );
OAI21X1 OAI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1565_), .B(_1507__bF_buf4), .C(_1566_), .Y(_341_) );
INVX2 INVX2_95 ( .gnd(gnd), .vdd(vdd), .A(regs_19__30_), .Y(_1567_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(wdata[30]), .B(_1507__bF_buf3), .Y(_1568_) );
OAI21X1 OAI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1567_), .B(_1507__bF_buf2), .C(_1568_), .Y(_343_) );
INVX2 INVX2_96 ( .gnd(gnd), .vdd(vdd), .A(regs_19__31_), .Y(_1569_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(wdata[31]), .B(_1507__bF_buf1), .Y(_1570_) );
OAI21X1 OAI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1569_), .B(_1507__bF_buf0), .C(_1570_), .Y(_344_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf8), .B(_1506__bF_buf4), .Y(_1571_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(regs_18__0_), .B(_1571__bF_buf7), .Y(_1572_) );
AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_992__bF_buf1), .B(_1571__bF_buf6), .C(_1572_), .Y(_288_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(regs_18__1_), .B(_1571__bF_buf5), .Y(_1573_) );
AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1003__bF_buf1), .B(_1571__bF_buf4), .C(_1573_), .Y(_299_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(regs_18__2_), .B(_1571__bF_buf3), .Y(_1574_) );
AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf1), .B(_1571__bF_buf2), .C(_1574_), .Y(_310_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(regs_18__3_), .B(_1571__bF_buf1), .Y(_1575_) );
AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1007__bF_buf1), .B(_1571__bF_buf0), .C(_1575_), .Y(_313_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(regs_18__4_), .B(_1571__bF_buf7), .Y(_1576_) );
AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1009__bF_buf0), .B(_1571__bF_buf6), .C(_1576_), .Y(_314_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(regs_18__5_), .B(_1571__bF_buf5), .Y(_1577_) );
AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1011__bF_buf0), .B(_1571__bF_buf4), .C(_1577_), .Y(_315_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(regs_18__6_), .B(_1571__bF_buf3), .Y(_1578_) );
AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1013__bF_buf0), .B(_1571__bF_buf2), .C(_1578_), .Y(_316_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(regs_18__7_), .B(_1571__bF_buf1), .Y(_1579_) );
AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1015__bF_buf0), .B(_1571__bF_buf0), .C(_1579_), .Y(_317_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(regs_18__8_), .B(_1571__bF_buf7), .Y(_1580_) );
AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf0), .B(_1571__bF_buf6), .C(_1580_), .Y(_318_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(regs_18__9_), .B(_1571__bF_buf5), .Y(_1581_) );
AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1019__bF_buf0), .B(_1571__bF_buf4), .C(_1581_), .Y(_319_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(regs_18__10_), .B(_1571__bF_buf3), .Y(_1582_) );
AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_1021__bF_buf0), .B(_1571__bF_buf2), .C(_1582_), .Y(_289_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(regs_18__11_), .B(_1571__bF_buf1), .Y(_1583_) );
AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_1023__bF_buf0), .B(_1571__bF_buf0), .C(_1583_), .Y(_290_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(regs_18__12_), .B(_1571__bF_buf7), .Y(_1584_) );
AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_1025__bF_buf0), .B(_1571__bF_buf6), .C(_1584_), .Y(_291_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(regs_18__13_), .B(_1571__bF_buf5), .Y(_1585_) );
AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_1027__bF_buf0), .B(_1571__bF_buf4), .C(_1585_), .Y(_292_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(regs_18__14_), .B(_1571__bF_buf3), .Y(_1586_) );
AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_1029__bF_buf0), .B(_1571__bF_buf2), .C(_1586_), .Y(_293_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(regs_18__15_), .B(_1571__bF_buf1), .Y(_1587_) );
AOI21X1 AOI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf0), .B(_1571__bF_buf0), .C(_1587_), .Y(_294_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(regs_18__16_), .B(_1571__bF_buf7), .Y(_1588_) );
AOI21X1 AOI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_1033__bF_buf0), .B(_1571__bF_buf6), .C(_1588_), .Y(_295_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(regs_18__17_), .B(_1571__bF_buf5), .Y(_1589_) );
AOI21X1 AOI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_1035__bF_buf0), .B(_1571__bF_buf4), .C(_1589_), .Y(_296_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(regs_18__18_), .B(_1571__bF_buf3), .Y(_1590_) );
AOI21X1 AOI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_1037__bF_buf0), .B(_1571__bF_buf2), .C(_1590_), .Y(_297_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(regs_18__19_), .B(_1571__bF_buf1), .Y(_1591_) );
AOI21X1 AOI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_1039__bF_buf0), .B(_1571__bF_buf0), .C(_1591_), .Y(_298_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(regs_18__20_), .B(_1571__bF_buf7), .Y(_1592_) );
AOI21X1 AOI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_1041__bF_buf0), .B(_1571__bF_buf6), .C(_1592_), .Y(_300_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(regs_18__21_), .B(_1571__bF_buf5), .Y(_1593_) );
AOI21X1 AOI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_1043__bF_buf0), .B(_1571__bF_buf4), .C(_1593_), .Y(_301_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(regs_18__22_), .B(_1571__bF_buf3), .Y(_1594_) );
AOI21X1 AOI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1045__bF_buf0), .B(_1571__bF_buf2), .C(_1594_), .Y(_302_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(regs_18__23_), .B(_1571__bF_buf1), .Y(_1595_) );
AOI21X1 AOI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_1047__bF_buf0), .B(_1571__bF_buf0), .C(_1595_), .Y(_303_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(regs_18__24_), .B(_1571__bF_buf7), .Y(_1596_) );
AOI21X1 AOI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1049__bF_buf0), .B(_1571__bF_buf6), .C(_1596_), .Y(_304_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(regs_18__25_), .B(_1571__bF_buf5), .Y(_1597_) );
AOI21X1 AOI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1051__bF_buf0), .B(_1571__bF_buf4), .C(_1597_), .Y(_305_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(regs_18__26_), .B(_1571__bF_buf3), .Y(_1598_) );
AOI21X1 AOI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_1053__bF_buf0), .B(_1571__bF_buf2), .C(_1598_), .Y(_306_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(regs_18__27_), .B(_1571__bF_buf1), .Y(_1599_) );
AOI21X1 AOI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_1055__bF_buf0), .B(_1571__bF_buf0), .C(_1599_), .Y(_307_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(regs_18__28_), .B(_1571__bF_buf7), .Y(_1600_) );
AOI21X1 AOI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_1057__bF_buf0), .B(_1571__bF_buf6), .C(_1600_), .Y(_308_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(regs_18__29_), .B(_1571__bF_buf5), .Y(_1601_) );
AOI21X1 AOI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_1059__bF_buf0), .B(_1571__bF_buf4), .C(_1601_), .Y(_309_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(regs_18__30_), .B(_1571__bF_buf3), .Y(_1602_) );
AOI21X1 AOI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_1061__bF_buf0), .B(_1571__bF_buf2), .C(_1602_), .Y(_311_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(regs_18__31_), .B(_1571__bF_buf1), .Y(_1603_) );
AOI21X1 AOI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_1063__bF_buf0), .B(_1571__bF_buf0), .C(_1603_), .Y(_312_) );
INVX2 INVX2_97 ( .gnd(gnd), .vdd(vdd), .A(regs_17__0_), .Y(_1604_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf3), .B(_1070__bF_buf9), .Y(_1605_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(wdata[0]), .B(_1605__bF_buf7), .Y(_1606_) );
OAI21X1 OAI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1604_), .B(_1605__bF_buf6), .C(_1606_), .Y(_256_) );
INVX2 INVX2_98 ( .gnd(gnd), .vdd(vdd), .A(regs_17__1_), .Y(_1607_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(wdata[1]), .B(_1605__bF_buf5), .Y(_1608_) );
OAI21X1 OAI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1607_), .B(_1605__bF_buf4), .C(_1608_), .Y(_267_) );
INVX2 INVX2_99 ( .gnd(gnd), .vdd(vdd), .A(regs_17__2_), .Y(_1609_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(wdata[2]), .B(_1605__bF_buf3), .Y(_1610_) );
OAI21X1 OAI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1609_), .B(_1605__bF_buf2), .C(_1610_), .Y(_278_) );
INVX2 INVX2_100 ( .gnd(gnd), .vdd(vdd), .A(regs_17__3_), .Y(_1611_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(wdata[3]), .B(_1605__bF_buf1), .Y(_1612_) );
OAI21X1 OAI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1611_), .B(_1605__bF_buf0), .C(_1612_), .Y(_281_) );
INVX2 INVX2_101 ( .gnd(gnd), .vdd(vdd), .A(regs_17__4_), .Y(_1613_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(wdata[4]), .B(_1605__bF_buf7), .Y(_1614_) );
OAI21X1 OAI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1613_), .B(_1605__bF_buf6), .C(_1614_), .Y(_282_) );
INVX2 INVX2_102 ( .gnd(gnd), .vdd(vdd), .A(regs_17__5_), .Y(_1615_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(wdata[5]), .B(_1605__bF_buf5), .Y(_1616_) );
OAI21X1 OAI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(_1605__bF_buf4), .C(_1616_), .Y(_283_) );
INVX2 INVX2_103 ( .gnd(gnd), .vdd(vdd), .A(regs_17__6_), .Y(_1617_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(wdata[6]), .B(_1605__bF_buf3), .Y(_1618_) );
OAI21X1 OAI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1617_), .B(_1605__bF_buf2), .C(_1618_), .Y(_284_) );
INVX2 INVX2_104 ( .gnd(gnd), .vdd(vdd), .A(regs_17__7_), .Y(_1619_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(wdata[7]), .B(_1605__bF_buf1), .Y(_1620_) );
OAI21X1 OAI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1619_), .B(_1605__bF_buf0), .C(_1620_), .Y(_285_) );
INVX2 INVX2_105 ( .gnd(gnd), .vdd(vdd), .A(regs_17__8_), .Y(_1621_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(wdata[8]), .B(_1605__bF_buf7), .Y(_1622_) );
OAI21X1 OAI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .B(_1605__bF_buf6), .C(_1622_), .Y(_286_) );
INVX2 INVX2_106 ( .gnd(gnd), .vdd(vdd), .A(regs_17__9_), .Y(_1623_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(wdata[9]), .B(_1605__bF_buf5), .Y(_1624_) );
OAI21X1 OAI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(_1605__bF_buf4), .C(_1624_), .Y(_287_) );
INVX2 INVX2_107 ( .gnd(gnd), .vdd(vdd), .A(regs_17__10_), .Y(_1625_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(wdata[10]), .B(_1605__bF_buf3), .Y(_1626_) );
OAI21X1 OAI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1625_), .B(_1605__bF_buf2), .C(_1626_), .Y(_257_) );
INVX2 INVX2_108 ( .gnd(gnd), .vdd(vdd), .A(regs_17__11_), .Y(_1627_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(wdata[11]), .B(_1605__bF_buf1), .Y(_1628_) );
OAI21X1 OAI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1627_), .B(_1605__bF_buf0), .C(_1628_), .Y(_258_) );
INVX2 INVX2_109 ( .gnd(gnd), .vdd(vdd), .A(regs_17__12_), .Y(_1629_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(wdata[12]), .B(_1605__bF_buf7), .Y(_1630_) );
OAI21X1 OAI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1629_), .B(_1605__bF_buf6), .C(_1630_), .Y(_259_) );
INVX2 INVX2_110 ( .gnd(gnd), .vdd(vdd), .A(regs_17__13_), .Y(_1631_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(wdata[13]), .B(_1605__bF_buf5), .Y(_1632_) );
OAI21X1 OAI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .B(_1605__bF_buf4), .C(_1632_), .Y(_260_) );
INVX2 INVX2_111 ( .gnd(gnd), .vdd(vdd), .A(regs_17__14_), .Y(_1633_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(wdata[14]), .B(_1605__bF_buf3), .Y(_1634_) );
OAI21X1 OAI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1633_), .B(_1605__bF_buf2), .C(_1634_), .Y(_261_) );
INVX2 INVX2_112 ( .gnd(gnd), .vdd(vdd), .A(regs_17__15_), .Y(_1635_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(wdata[15]), .B(_1605__bF_buf1), .Y(_1636_) );
OAI21X1 OAI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .B(_1605__bF_buf0), .C(_1636_), .Y(_262_) );
INVX2 INVX2_113 ( .gnd(gnd), .vdd(vdd), .A(regs_17__16_), .Y(_1637_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(wdata[16]), .B(_1605__bF_buf7), .Y(_1638_) );
OAI21X1 OAI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1637_), .B(_1605__bF_buf6), .C(_1638_), .Y(_263_) );
INVX2 INVX2_114 ( .gnd(gnd), .vdd(vdd), .A(regs_17__17_), .Y(_1639_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(wdata[17]), .B(_1605__bF_buf5), .Y(_1640_) );
OAI21X1 OAI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .B(_1605__bF_buf4), .C(_1640_), .Y(_264_) );
INVX2 INVX2_115 ( .gnd(gnd), .vdd(vdd), .A(regs_17__18_), .Y(_1641_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(wdata[18]), .B(_1605__bF_buf3), .Y(_1642_) );
OAI21X1 OAI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1641_), .B(_1605__bF_buf2), .C(_1642_), .Y(_265_) );
INVX2 INVX2_116 ( .gnd(gnd), .vdd(vdd), .A(regs_17__19_), .Y(_1643_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(wdata[19]), .B(_1605__bF_buf1), .Y(_1644_) );
OAI21X1 OAI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .B(_1605__bF_buf0), .C(_1644_), .Y(_266_) );
INVX2 INVX2_117 ( .gnd(gnd), .vdd(vdd), .A(regs_17__20_), .Y(_1645_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(wdata[20]), .B(_1605__bF_buf7), .Y(_1646_) );
OAI21X1 OAI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1645_), .B(_1605__bF_buf6), .C(_1646_), .Y(_268_) );
INVX2 INVX2_118 ( .gnd(gnd), .vdd(vdd), .A(regs_17__21_), .Y(_1647_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(wdata[21]), .B(_1605__bF_buf5), .Y(_1648_) );
OAI21X1 OAI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1647_), .B(_1605__bF_buf4), .C(_1648_), .Y(_269_) );
INVX2 INVX2_119 ( .gnd(gnd), .vdd(vdd), .A(regs_17__22_), .Y(_1649_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(wdata[22]), .B(_1605__bF_buf3), .Y(_1650_) );
OAI21X1 OAI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1649_), .B(_1605__bF_buf2), .C(_1650_), .Y(_270_) );
INVX2 INVX2_120 ( .gnd(gnd), .vdd(vdd), .A(regs_17__23_), .Y(_1651_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(wdata[23]), .B(_1605__bF_buf1), .Y(_1652_) );
OAI21X1 OAI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1651_), .B(_1605__bF_buf0), .C(_1652_), .Y(_271_) );
INVX2 INVX2_121 ( .gnd(gnd), .vdd(vdd), .A(regs_17__24_), .Y(_1653_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(wdata[24]), .B(_1605__bF_buf7), .Y(_1654_) );
OAI21X1 OAI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .B(_1605__bF_buf6), .C(_1654_), .Y(_272_) );
INVX2 INVX2_122 ( .gnd(gnd), .vdd(vdd), .A(regs_17__25_), .Y(_1655_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(wdata[25]), .B(_1605__bF_buf5), .Y(_1656_) );
OAI21X1 OAI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .B(_1605__bF_buf4), .C(_1656_), .Y(_273_) );
INVX2 INVX2_123 ( .gnd(gnd), .vdd(vdd), .A(regs_17__26_), .Y(_1657_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(wdata[26]), .B(_1605__bF_buf3), .Y(_1658_) );
OAI21X1 OAI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1657_), .B(_1605__bF_buf2), .C(_1658_), .Y(_274_) );
INVX2 INVX2_124 ( .gnd(gnd), .vdd(vdd), .A(regs_17__27_), .Y(_1659_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(wdata[27]), .B(_1605__bF_buf1), .Y(_1660_) );
OAI21X1 OAI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_1659_), .B(_1605__bF_buf0), .C(_1660_), .Y(_275_) );
INVX2 INVX2_125 ( .gnd(gnd), .vdd(vdd), .A(regs_17__28_), .Y(_1661_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(wdata[28]), .B(_1605__bF_buf7), .Y(_1662_) );
OAI21X1 OAI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1661_), .B(_1605__bF_buf6), .C(_1662_), .Y(_276_) );
INVX2 INVX2_126 ( .gnd(gnd), .vdd(vdd), .A(regs_17__29_), .Y(_1663_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(wdata[29]), .B(_1605__bF_buf5), .Y(_1664_) );
OAI21X1 OAI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1663_), .B(_1605__bF_buf4), .C(_1664_), .Y(_277_) );
INVX2 INVX2_127 ( .gnd(gnd), .vdd(vdd), .A(regs_17__30_), .Y(_1665_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(wdata[30]), .B(_1605__bF_buf3), .Y(_1666_) );
OAI21X1 OAI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_1665_), .B(_1605__bF_buf2), .C(_1666_), .Y(_279_) );
INVX2 INVX2_128 ( .gnd(gnd), .vdd(vdd), .A(regs_17__31_), .Y(_1667_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(wdata[31]), .B(_1605__bF_buf1), .Y(_1668_) );
OAI21X1 OAI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1667_), .B(_1605__bF_buf0), .C(_1668_), .Y(_280_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf2), .B(_1104__bF_buf13), .Y(_1669_) );
OAI21X1 OAI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf1), .B(_1104__bF_buf12), .C(regs_16__0_), .Y(_1670_) );
OAI21X1 OAI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf4), .B(_992__bF_buf0), .C(_1670_), .Y(_224_) );
OAI21X1 OAI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf0), .B(_1104__bF_buf11), .C(regs_16__1_), .Y(_1671_) );
OAI21X1 OAI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf3), .B(_1003__bF_buf0), .C(_1671_), .Y(_235_) );
OAI21X1 OAI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf5), .B(_1104__bF_buf10), .C(regs_16__2_), .Y(_1672_) );
OAI21X1 OAI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf2), .B(_1005__bF_buf0), .C(_1672_), .Y(_246_) );
OAI21X1 OAI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf4), .B(_1104__bF_buf9), .C(regs_16__3_), .Y(_1673_) );
OAI21X1 OAI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf1), .B(_1007__bF_buf0), .C(_1673_), .Y(_249_) );
OAI21X1 OAI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf3), .B(_1104__bF_buf8), .C(regs_16__4_), .Y(_1674_) );
OAI21X1 OAI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf0), .B(_1009__bF_buf3), .C(_1674_), .Y(_250_) );
OAI21X1 OAI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf2), .B(_1104__bF_buf7), .C(regs_16__5_), .Y(_1675_) );
OAI21X1 OAI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf4), .B(_1011__bF_buf3), .C(_1675_), .Y(_251_) );
OAI21X1 OAI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf1), .B(_1104__bF_buf6), .C(regs_16__6_), .Y(_1676_) );
OAI21X1 OAI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf3), .B(_1013__bF_buf3), .C(_1676_), .Y(_252_) );
OAI21X1 OAI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf0), .B(_1104__bF_buf5), .C(regs_16__7_), .Y(_1677_) );
OAI21X1 OAI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf2), .B(_1015__bF_buf3), .C(_1677_), .Y(_253_) );
OAI21X1 OAI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf5), .B(_1104__bF_buf4), .C(regs_16__8_), .Y(_1678_) );
OAI21X1 OAI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf1), .B(_1017__bF_buf3), .C(_1678_), .Y(_254_) );
OAI21X1 OAI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf4), .B(_1104__bF_buf3), .C(regs_16__9_), .Y(_1679_) );
OAI21X1 OAI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf0), .B(_1019__bF_buf3), .C(_1679_), .Y(_255_) );
OAI21X1 OAI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf3), .B(_1104__bF_buf2), .C(regs_16__10_), .Y(_1680_) );
OAI21X1 OAI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf4), .B(_1021__bF_buf3), .C(_1680_), .Y(_225_) );
OAI21X1 OAI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf2), .B(_1104__bF_buf1), .C(regs_16__11_), .Y(_1681_) );
OAI21X1 OAI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf3), .B(_1023__bF_buf3), .C(_1681_), .Y(_226_) );
OAI21X1 OAI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf1), .B(_1104__bF_buf0), .C(regs_16__12_), .Y(_1682_) );
OAI21X1 OAI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf2), .B(_1025__bF_buf3), .C(_1682_), .Y(_227_) );
OAI21X1 OAI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf0), .B(_1104__bF_buf14), .C(regs_16__13_), .Y(_1683_) );
OAI21X1 OAI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf1), .B(_1027__bF_buf3), .C(_1683_), .Y(_228_) );
OAI21X1 OAI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf5), .B(_1104__bF_buf13), .C(regs_16__14_), .Y(_1684_) );
OAI21X1 OAI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf0), .B(_1029__bF_buf3), .C(_1684_), .Y(_229_) );
OAI21X1 OAI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf4), .B(_1104__bF_buf12), .C(regs_16__15_), .Y(_1685_) );
OAI21X1 OAI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf4), .B(_1031__bF_buf3), .C(_1685_), .Y(_230_) );
OAI21X1 OAI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf3), .B(_1104__bF_buf11), .C(regs_16__16_), .Y(_1686_) );
OAI21X1 OAI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf3), .B(_1033__bF_buf3), .C(_1686_), .Y(_231_) );
OAI21X1 OAI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf2), .B(_1104__bF_buf10), .C(regs_16__17_), .Y(_1687_) );
OAI21X1 OAI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf2), .B(_1035__bF_buf3), .C(_1687_), .Y(_232_) );
OAI21X1 OAI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf1), .B(_1104__bF_buf9), .C(regs_16__18_), .Y(_1688_) );
OAI21X1 OAI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf1), .B(_1037__bF_buf3), .C(_1688_), .Y(_233_) );
OAI21X1 OAI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf0), .B(_1104__bF_buf8), .C(regs_16__19_), .Y(_1689_) );
OAI21X1 OAI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf0), .B(_1039__bF_buf3), .C(_1689_), .Y(_234_) );
OAI21X1 OAI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf5), .B(_1104__bF_buf7), .C(regs_16__20_), .Y(_1690_) );
OAI21X1 OAI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf4), .B(_1041__bF_buf3), .C(_1690_), .Y(_236_) );
OAI21X1 OAI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf4), .B(_1104__bF_buf6), .C(regs_16__21_), .Y(_1691_) );
OAI21X1 OAI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf3), .B(_1043__bF_buf3), .C(_1691_), .Y(_237_) );
OAI21X1 OAI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf3), .B(_1104__bF_buf5), .C(regs_16__22_), .Y(_1692_) );
OAI21X1 OAI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf2), .B(_1045__bF_buf3), .C(_1692_), .Y(_238_) );
OAI21X1 OAI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf2), .B(_1104__bF_buf4), .C(regs_16__23_), .Y(_1693_) );
OAI21X1 OAI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf1), .B(_1047__bF_buf3), .C(_1693_), .Y(_239_) );
OAI21X1 OAI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf1), .B(_1104__bF_buf3), .C(regs_16__24_), .Y(_1694_) );
OAI21X1 OAI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf0), .B(_1049__bF_buf3), .C(_1694_), .Y(_240_) );
OAI21X1 OAI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf0), .B(_1104__bF_buf2), .C(regs_16__25_), .Y(_1695_) );
OAI21X1 OAI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf4), .B(_1051__bF_buf3), .C(_1695_), .Y(_241_) );
OAI21X1 OAI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf5), .B(_1104__bF_buf1), .C(regs_16__26_), .Y(_1696_) );
OAI21X1 OAI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf3), .B(_1053__bF_buf3), .C(_1696_), .Y(_242_) );
OAI21X1 OAI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf4), .B(_1104__bF_buf0), .C(regs_16__27_), .Y(_1697_) );
OAI21X1 OAI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf2), .B(_1055__bF_buf3), .C(_1697_), .Y(_243_) );
OAI21X1 OAI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf3), .B(_1104__bF_buf14), .C(regs_16__28_), .Y(_1698_) );
OAI21X1 OAI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf1), .B(_1057__bF_buf3), .C(_1698_), .Y(_244_) );
OAI21X1 OAI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf2), .B(_1104__bF_buf13), .C(regs_16__29_), .Y(_1699_) );
OAI21X1 OAI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf0), .B(_1059__bF_buf3), .C(_1699_), .Y(_245_) );
OAI21X1 OAI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf1), .B(_1104__bF_buf12), .C(regs_16__30_), .Y(_1700_) );
OAI21X1 OAI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf4), .B(_1061__bF_buf3), .C(_1700_), .Y(_247_) );
OAI21X1 OAI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_1506__bF_buf0), .B(_1104__bF_buf11), .C(regs_16__31_), .Y(_1701_) );
OAI21X1 OAI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_1669__bF_buf3), .B(_1063__bF_buf3), .C(_1701_), .Y(_248_) );
INVX2 INVX2_129 ( .gnd(gnd), .vdd(vdd), .A(regs_15__0_), .Y(_1702_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(waddr[4]), .B(_994_), .Y(_1703_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_1703_), .B(waddr[2]), .Y(_1704_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1142__bF_buf3), .B(_1704__bF_buf5), .Y(_1705_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(wdata[0]), .B(_1705__bF_buf7), .Y(_1706_) );
OAI21X1 OAI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(_1702_), .B(_1705__bF_buf6), .C(_1706_), .Y(_192_) );
INVX2 INVX2_130 ( .gnd(gnd), .vdd(vdd), .A(regs_15__1_), .Y(_1707_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(wdata[1]), .B(_1705__bF_buf5), .Y(_1708_) );
OAI21X1 OAI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_1707_), .B(_1705__bF_buf4), .C(_1708_), .Y(_203_) );
INVX2 INVX2_131 ( .gnd(gnd), .vdd(vdd), .A(regs_15__2_), .Y(_1709_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(wdata[2]), .B(_1705__bF_buf3), .Y(_1710_) );
OAI21X1 OAI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_1709_), .B(_1705__bF_buf2), .C(_1710_), .Y(_214_) );
INVX2 INVX2_132 ( .gnd(gnd), .vdd(vdd), .A(regs_15__3_), .Y(_1711_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(wdata[3]), .B(_1705__bF_buf1), .Y(_1712_) );
OAI21X1 OAI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_1711_), .B(_1705__bF_buf0), .C(_1712_), .Y(_217_) );
INVX2 INVX2_133 ( .gnd(gnd), .vdd(vdd), .A(regs_15__4_), .Y(_1713_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(wdata[4]), .B(_1705__bF_buf7), .Y(_1714_) );
OAI21X1 OAI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_1713_), .B(_1705__bF_buf6), .C(_1714_), .Y(_218_) );
INVX2 INVX2_134 ( .gnd(gnd), .vdd(vdd), .A(regs_15__5_), .Y(_1715_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(wdata[5]), .B(_1705__bF_buf5), .Y(_1716_) );
OAI21X1 OAI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(_1715_), .B(_1705__bF_buf4), .C(_1716_), .Y(_219_) );
INVX2 INVX2_135 ( .gnd(gnd), .vdd(vdd), .A(regs_15__6_), .Y(_1717_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(wdata[6]), .B(_1705__bF_buf3), .Y(_1718_) );
OAI21X1 OAI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(_1717_), .B(_1705__bF_buf2), .C(_1718_), .Y(_220_) );
INVX2 INVX2_136 ( .gnd(gnd), .vdd(vdd), .A(regs_15__7_), .Y(_1719_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(wdata[7]), .B(_1705__bF_buf1), .Y(_1720_) );
OAI21X1 OAI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_1719_), .B(_1705__bF_buf0), .C(_1720_), .Y(_221_) );
INVX2 INVX2_137 ( .gnd(gnd), .vdd(vdd), .A(regs_15__8_), .Y(_1721_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(wdata[8]), .B(_1705__bF_buf7), .Y(_1722_) );
OAI21X1 OAI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_1721_), .B(_1705__bF_buf6), .C(_1722_), .Y(_222_) );
INVX2 INVX2_138 ( .gnd(gnd), .vdd(vdd), .A(regs_15__9_), .Y(_1723_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(wdata[9]), .B(_1705__bF_buf5), .Y(_1724_) );
OAI21X1 OAI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_1723_), .B(_1705__bF_buf4), .C(_1724_), .Y(_223_) );
INVX2 INVX2_139 ( .gnd(gnd), .vdd(vdd), .A(regs_15__10_), .Y(_1725_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(wdata[10]), .B(_1705__bF_buf3), .Y(_1726_) );
OAI21X1 OAI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_1725_), .B(_1705__bF_buf2), .C(_1726_), .Y(_193_) );
INVX2 INVX2_140 ( .gnd(gnd), .vdd(vdd), .A(regs_15__11_), .Y(_1727_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(wdata[11]), .B(_1705__bF_buf1), .Y(_1728_) );
OAI21X1 OAI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(_1727_), .B(_1705__bF_buf0), .C(_1728_), .Y(_194_) );
INVX2 INVX2_141 ( .gnd(gnd), .vdd(vdd), .A(regs_15__12_), .Y(_1729_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(wdata[12]), .B(_1705__bF_buf7), .Y(_1730_) );
OAI21X1 OAI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(_1729_), .B(_1705__bF_buf6), .C(_1730_), .Y(_195_) );
INVX2 INVX2_142 ( .gnd(gnd), .vdd(vdd), .A(regs_15__13_), .Y(_1731_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(wdata[13]), .B(_1705__bF_buf5), .Y(_1732_) );
OAI21X1 OAI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_1731_), .B(_1705__bF_buf4), .C(_1732_), .Y(_196_) );
INVX2 INVX2_143 ( .gnd(gnd), .vdd(vdd), .A(regs_15__14_), .Y(_1733_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(wdata[14]), .B(_1705__bF_buf3), .Y(_1734_) );
OAI21X1 OAI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(_1733_), .B(_1705__bF_buf2), .C(_1734_), .Y(_197_) );
INVX2 INVX2_144 ( .gnd(gnd), .vdd(vdd), .A(regs_15__15_), .Y(_1735_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(wdata[15]), .B(_1705__bF_buf1), .Y(_1736_) );
OAI21X1 OAI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .B(_1705__bF_buf0), .C(_1736_), .Y(_198_) );
INVX2 INVX2_145 ( .gnd(gnd), .vdd(vdd), .A(regs_15__16_), .Y(_1737_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(wdata[16]), .B(_1705__bF_buf7), .Y(_1738_) );
OAI21X1 OAI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1705__bF_buf6), .C(_1738_), .Y(_199_) );
INVX2 INVX2_146 ( .gnd(gnd), .vdd(vdd), .A(regs_15__17_), .Y(_1739_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(wdata[17]), .B(_1705__bF_buf5), .Y(_1740_) );
OAI21X1 OAI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(_1739_), .B(_1705__bF_buf4), .C(_1740_), .Y(_200_) );
INVX2 INVX2_147 ( .gnd(gnd), .vdd(vdd), .A(regs_15__18_), .Y(_1741_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(wdata[18]), .B(_1705__bF_buf3), .Y(_1742_) );
OAI21X1 OAI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_1741_), .B(_1705__bF_buf2), .C(_1742_), .Y(_201_) );
INVX2 INVX2_148 ( .gnd(gnd), .vdd(vdd), .A(regs_15__19_), .Y(_1743_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(wdata[19]), .B(_1705__bF_buf1), .Y(_1744_) );
OAI21X1 OAI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_1743_), .B(_1705__bF_buf0), .C(_1744_), .Y(_202_) );
INVX2 INVX2_149 ( .gnd(gnd), .vdd(vdd), .A(regs_15__20_), .Y(_1745_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(wdata[20]), .B(_1705__bF_buf7), .Y(_1746_) );
OAI21X1 OAI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(_1745_), .B(_1705__bF_buf6), .C(_1746_), .Y(_204_) );
INVX2 INVX2_150 ( .gnd(gnd), .vdd(vdd), .A(regs_15__21_), .Y(_1747_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(wdata[21]), .B(_1705__bF_buf5), .Y(_1748_) );
OAI21X1 OAI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_1747_), .B(_1705__bF_buf4), .C(_1748_), .Y(_205_) );
INVX2 INVX2_151 ( .gnd(gnd), .vdd(vdd), .A(regs_15__22_), .Y(_1749_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(wdata[22]), .B(_1705__bF_buf3), .Y(_1750_) );
OAI21X1 OAI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_1749_), .B(_1705__bF_buf2), .C(_1750_), .Y(_206_) );
INVX2 INVX2_152 ( .gnd(gnd), .vdd(vdd), .A(regs_15__23_), .Y(_1751_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(wdata[23]), .B(_1705__bF_buf1), .Y(_1752_) );
OAI21X1 OAI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_1751_), .B(_1705__bF_buf0), .C(_1752_), .Y(_207_) );
INVX2 INVX2_153 ( .gnd(gnd), .vdd(vdd), .A(regs_15__24_), .Y(_1753_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(wdata[24]), .B(_1705__bF_buf7), .Y(_1754_) );
OAI21X1 OAI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(_1753_), .B(_1705__bF_buf6), .C(_1754_), .Y(_208_) );
INVX2 INVX2_154 ( .gnd(gnd), .vdd(vdd), .A(regs_15__25_), .Y(_1755_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(wdata[25]), .B(_1705__bF_buf5), .Y(_1756_) );
OAI21X1 OAI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(_1755_), .B(_1705__bF_buf4), .C(_1756_), .Y(_209_) );
INVX2 INVX2_155 ( .gnd(gnd), .vdd(vdd), .A(regs_15__26_), .Y(_1757_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(wdata[26]), .B(_1705__bF_buf3), .Y(_1758_) );
OAI21X1 OAI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_1757_), .B(_1705__bF_buf2), .C(_1758_), .Y(_210_) );
INVX2 INVX2_156 ( .gnd(gnd), .vdd(vdd), .A(regs_15__27_), .Y(_1759_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(wdata[27]), .B(_1705__bF_buf1), .Y(_1760_) );
OAI21X1 OAI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(_1759_), .B(_1705__bF_buf0), .C(_1760_), .Y(_211_) );
INVX2 INVX2_157 ( .gnd(gnd), .vdd(vdd), .A(regs_15__28_), .Y(_1761_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(wdata[28]), .B(_1705__bF_buf7), .Y(_1762_) );
OAI21X1 OAI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_1761_), .B(_1705__bF_buf6), .C(_1762_), .Y(_212_) );
INVX2 INVX2_158 ( .gnd(gnd), .vdd(vdd), .A(regs_15__29_), .Y(_1763_) );
NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(wdata[29]), .B(_1705__bF_buf5), .Y(_1764_) );
OAI21X1 OAI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_1763_), .B(_1705__bF_buf4), .C(_1764_), .Y(_213_) );
INVX2 INVX2_159 ( .gnd(gnd), .vdd(vdd), .A(regs_15__30_), .Y(_1765_) );
NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(wdata[30]), .B(_1705__bF_buf3), .Y(_1766_) );
OAI21X1 OAI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_1765_), .B(_1705__bF_buf2), .C(_1766_), .Y(_215_) );
INVX2 INVX2_160 ( .gnd(gnd), .vdd(vdd), .A(regs_15__31_), .Y(_1767_) );
NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(wdata[31]), .B(_1705__bF_buf1), .Y(_1768_) );
OAI21X1 OAI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(_1767_), .B(_1705__bF_buf0), .C(_1768_), .Y(_216_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf7), .B(_1704__bF_buf4), .Y(_1769_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(regs_14__0_), .B(_1769__bF_buf7), .Y(_1770_) );
AOI21X1 AOI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_992__bF_buf3), .B(_1769__bF_buf6), .C(_1770_), .Y(_160_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(regs_14__1_), .B(_1769__bF_buf5), .Y(_1771_) );
AOI21X1 AOI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_1003__bF_buf3), .B(_1769__bF_buf4), .C(_1771_), .Y(_171_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(regs_14__2_), .B(_1769__bF_buf3), .Y(_1772_) );
AOI21X1 AOI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf3), .B(_1769__bF_buf2), .C(_1772_), .Y(_182_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(regs_14__3_), .B(_1769__bF_buf1), .Y(_1773_) );
AOI21X1 AOI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_1007__bF_buf3), .B(_1769__bF_buf0), .C(_1773_), .Y(_185_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(regs_14__4_), .B(_1769__bF_buf7), .Y(_1774_) );
AOI21X1 AOI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_1009__bF_buf2), .B(_1769__bF_buf6), .C(_1774_), .Y(_186_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(regs_14__5_), .B(_1769__bF_buf5), .Y(_1775_) );
AOI21X1 AOI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_1011__bF_buf2), .B(_1769__bF_buf4), .C(_1775_), .Y(_187_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(regs_14__6_), .B(_1769__bF_buf3), .Y(_1776_) );
AOI21X1 AOI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_1013__bF_buf2), .B(_1769__bF_buf2), .C(_1776_), .Y(_188_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(regs_14__7_), .B(_1769__bF_buf1), .Y(_1777_) );
AOI21X1 AOI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_1015__bF_buf2), .B(_1769__bF_buf0), .C(_1777_), .Y(_189_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(regs_14__8_), .B(_1769__bF_buf7), .Y(_1778_) );
AOI21X1 AOI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf2), .B(_1769__bF_buf6), .C(_1778_), .Y(_190_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(regs_14__9_), .B(_1769__bF_buf5), .Y(_1779_) );
AOI21X1 AOI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_1019__bF_buf2), .B(_1769__bF_buf4), .C(_1779_), .Y(_191_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(regs_14__10_), .B(_1769__bF_buf3), .Y(_1780_) );
AOI21X1 AOI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_1021__bF_buf2), .B(_1769__bF_buf2), .C(_1780_), .Y(_161_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(regs_14__11_), .B(_1769__bF_buf1), .Y(_1781_) );
AOI21X1 AOI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_1023__bF_buf2), .B(_1769__bF_buf0), .C(_1781_), .Y(_162_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(regs_14__12_), .B(_1769__bF_buf7), .Y(_1782_) );
AOI21X1 AOI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_1025__bF_buf2), .B(_1769__bF_buf6), .C(_1782_), .Y(_163_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(regs_14__13_), .B(_1769__bF_buf5), .Y(_1783_) );
AOI21X1 AOI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1027__bF_buf2), .B(_1769__bF_buf4), .C(_1783_), .Y(_164_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(regs_14__14_), .B(_1769__bF_buf3), .Y(_1784_) );
AOI21X1 AOI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_1029__bF_buf2), .B(_1769__bF_buf2), .C(_1784_), .Y(_165_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(regs_14__15_), .B(_1769__bF_buf1), .Y(_1785_) );
AOI21X1 AOI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf2), .B(_1769__bF_buf0), .C(_1785_), .Y(_166_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(regs_14__16_), .B(_1769__bF_buf7), .Y(_1786_) );
AOI21X1 AOI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1033__bF_buf2), .B(_1769__bF_buf6), .C(_1786_), .Y(_167_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(regs_14__17_), .B(_1769__bF_buf5), .Y(_1787_) );
AOI21X1 AOI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1035__bF_buf2), .B(_1769__bF_buf4), .C(_1787_), .Y(_168_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(regs_14__18_), .B(_1769__bF_buf3), .Y(_1788_) );
AOI21X1 AOI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1037__bF_buf2), .B(_1769__bF_buf2), .C(_1788_), .Y(_169_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(regs_14__19_), .B(_1769__bF_buf1), .Y(_1789_) );
AOI21X1 AOI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_1039__bF_buf2), .B(_1769__bF_buf0), .C(_1789_), .Y(_170_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(regs_14__20_), .B(_1769__bF_buf7), .Y(_1790_) );
AOI21X1 AOI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1041__bF_buf2), .B(_1769__bF_buf6), .C(_1790_), .Y(_172_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(regs_14__21_), .B(_1769__bF_buf5), .Y(_1791_) );
AOI21X1 AOI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1043__bF_buf2), .B(_1769__bF_buf4), .C(_1791_), .Y(_173_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(regs_14__22_), .B(_1769__bF_buf3), .Y(_1792_) );
AOI21X1 AOI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1045__bF_buf2), .B(_1769__bF_buf2), .C(_1792_), .Y(_174_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(regs_14__23_), .B(_1769__bF_buf1), .Y(_1793_) );
AOI21X1 AOI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1047__bF_buf2), .B(_1769__bF_buf0), .C(_1793_), .Y(_175_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(regs_14__24_), .B(_1769__bF_buf7), .Y(_1794_) );
AOI21X1 AOI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1049__bF_buf2), .B(_1769__bF_buf6), .C(_1794_), .Y(_176_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(regs_14__25_), .B(_1769__bF_buf5), .Y(_1795_) );
AOI21X1 AOI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1051__bF_buf2), .B(_1769__bF_buf4), .C(_1795_), .Y(_177_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(regs_14__26_), .B(_1769__bF_buf3), .Y(_1796_) );
AOI21X1 AOI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1053__bF_buf2), .B(_1769__bF_buf2), .C(_1796_), .Y(_178_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(regs_14__27_), .B(_1769__bF_buf1), .Y(_1797_) );
AOI21X1 AOI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1055__bF_buf2), .B(_1769__bF_buf0), .C(_1797_), .Y(_179_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(regs_14__28_), .B(_1769__bF_buf7), .Y(_1798_) );
AOI21X1 AOI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_1057__bF_buf2), .B(_1769__bF_buf6), .C(_1798_), .Y(_180_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(regs_14__29_), .B(_1769__bF_buf5), .Y(_1799_) );
AOI21X1 AOI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1059__bF_buf2), .B(_1769__bF_buf4), .C(_1799_), .Y(_181_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(regs_14__30_), .B(_1769__bF_buf3), .Y(_1800_) );
AOI21X1 AOI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1061__bF_buf2), .B(_1769__bF_buf2), .C(_1800_), .Y(_183_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(regs_14__31_), .B(_1769__bF_buf1), .Y(_1801_) );
AOI21X1 AOI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1063__bF_buf2), .B(_1769__bF_buf0), .C(_1801_), .Y(_184_) );
INVX2 INVX2_161 ( .gnd(gnd), .vdd(vdd), .A(regs_13__0_), .Y(_1802_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf3), .B(_1070__bF_buf8), .Y(_1803_) );
NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(wdata[0]), .B(_1803__bF_buf7), .Y(_1804_) );
OAI21X1 OAI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_1802_), .B(_1803__bF_buf6), .C(_1804_), .Y(_128_) );
INVX2 INVX2_162 ( .gnd(gnd), .vdd(vdd), .A(regs_13__1_), .Y(_1805_) );
NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(wdata[1]), .B(_1803__bF_buf5), .Y(_1806_) );
OAI21X1 OAI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_1805_), .B(_1803__bF_buf4), .C(_1806_), .Y(_139_) );
INVX2 INVX2_163 ( .gnd(gnd), .vdd(vdd), .A(regs_13__2_), .Y(_1807_) );
NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(wdata[2]), .B(_1803__bF_buf3), .Y(_1808_) );
OAI21X1 OAI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_1807_), .B(_1803__bF_buf2), .C(_1808_), .Y(_150_) );
INVX2 INVX2_164 ( .gnd(gnd), .vdd(vdd), .A(regs_13__3_), .Y(_1809_) );
NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(wdata[3]), .B(_1803__bF_buf1), .Y(_1810_) );
OAI21X1 OAI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_1809_), .B(_1803__bF_buf0), .C(_1810_), .Y(_153_) );
INVX2 INVX2_165 ( .gnd(gnd), .vdd(vdd), .A(regs_13__4_), .Y(_1811_) );
NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(wdata[4]), .B(_1803__bF_buf7), .Y(_1812_) );
OAI21X1 OAI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_1811_), .B(_1803__bF_buf6), .C(_1812_), .Y(_154_) );
INVX2 INVX2_166 ( .gnd(gnd), .vdd(vdd), .A(regs_13__5_), .Y(_1813_) );
NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(wdata[5]), .B(_1803__bF_buf5), .Y(_1814_) );
OAI21X1 OAI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_1813_), .B(_1803__bF_buf4), .C(_1814_), .Y(_155_) );
INVX2 INVX2_167 ( .gnd(gnd), .vdd(vdd), .A(regs_13__6_), .Y(_1815_) );
NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(wdata[6]), .B(_1803__bF_buf3), .Y(_1816_) );
OAI21X1 OAI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_1815_), .B(_1803__bF_buf2), .C(_1816_), .Y(_156_) );
INVX2 INVX2_168 ( .gnd(gnd), .vdd(vdd), .A(regs_13__7_), .Y(_1817_) );
NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(wdata[7]), .B(_1803__bF_buf1), .Y(_1818_) );
OAI21X1 OAI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(_1817_), .B(_1803__bF_buf0), .C(_1818_), .Y(_157_) );
INVX2 INVX2_169 ( .gnd(gnd), .vdd(vdd), .A(regs_13__8_), .Y(_1819_) );
NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(wdata[8]), .B(_1803__bF_buf7), .Y(_1820_) );
OAI21X1 OAI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_1819_), .B(_1803__bF_buf6), .C(_1820_), .Y(_158_) );
INVX2 INVX2_170 ( .gnd(gnd), .vdd(vdd), .A(regs_13__9_), .Y(_1821_) );
NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(wdata[9]), .B(_1803__bF_buf5), .Y(_1822_) );
OAI21X1 OAI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_1821_), .B(_1803__bF_buf4), .C(_1822_), .Y(_159_) );
INVX2 INVX2_171 ( .gnd(gnd), .vdd(vdd), .A(regs_13__10_), .Y(_1823_) );
NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(wdata[10]), .B(_1803__bF_buf3), .Y(_1824_) );
OAI21X1 OAI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_1823_), .B(_1803__bF_buf2), .C(_1824_), .Y(_129_) );
INVX2 INVX2_172 ( .gnd(gnd), .vdd(vdd), .A(regs_13__11_), .Y(_1825_) );
NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(wdata[11]), .B(_1803__bF_buf1), .Y(_1826_) );
OAI21X1 OAI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_1825_), .B(_1803__bF_buf0), .C(_1826_), .Y(_130_) );
INVX2 INVX2_173 ( .gnd(gnd), .vdd(vdd), .A(regs_13__12_), .Y(_1827_) );
NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(wdata[12]), .B(_1803__bF_buf7), .Y(_1828_) );
OAI21X1 OAI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .B(_1803__bF_buf6), .C(_1828_), .Y(_131_) );
INVX2 INVX2_174 ( .gnd(gnd), .vdd(vdd), .A(regs_13__13_), .Y(_1829_) );
NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(wdata[13]), .B(_1803__bF_buf5), .Y(_1830_) );
OAI21X1 OAI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(_1829_), .B(_1803__bF_buf4), .C(_1830_), .Y(_132_) );
INVX2 INVX2_175 ( .gnd(gnd), .vdd(vdd), .A(regs_13__14_), .Y(_1831_) );
NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(wdata[14]), .B(_1803__bF_buf3), .Y(_1832_) );
OAI21X1 OAI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_1831_), .B(_1803__bF_buf2), .C(_1832_), .Y(_133_) );
INVX2 INVX2_176 ( .gnd(gnd), .vdd(vdd), .A(regs_13__15_), .Y(_1833_) );
NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(wdata[15]), .B(_1803__bF_buf1), .Y(_1834_) );
OAI21X1 OAI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_1833_), .B(_1803__bF_buf0), .C(_1834_), .Y(_134_) );
INVX2 INVX2_177 ( .gnd(gnd), .vdd(vdd), .A(regs_13__16_), .Y(_1835_) );
NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(wdata[16]), .B(_1803__bF_buf7), .Y(_1836_) );
OAI21X1 OAI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_1835_), .B(_1803__bF_buf6), .C(_1836_), .Y(_135_) );
INVX2 INVX2_178 ( .gnd(gnd), .vdd(vdd), .A(regs_13__17_), .Y(_1837_) );
NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(wdata[17]), .B(_1803__bF_buf5), .Y(_1838_) );
OAI21X1 OAI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_1837_), .B(_1803__bF_buf4), .C(_1838_), .Y(_136_) );
INVX2 INVX2_179 ( .gnd(gnd), .vdd(vdd), .A(regs_13__18_), .Y(_1839_) );
NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(wdata[18]), .B(_1803__bF_buf3), .Y(_1840_) );
OAI21X1 OAI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_1839_), .B(_1803__bF_buf2), .C(_1840_), .Y(_137_) );
INVX2 INVX2_180 ( .gnd(gnd), .vdd(vdd), .A(regs_13__19_), .Y(_1841_) );
NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(wdata[19]), .B(_1803__bF_buf1), .Y(_1842_) );
OAI21X1 OAI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_1841_), .B(_1803__bF_buf0), .C(_1842_), .Y(_138_) );
INVX2 INVX2_181 ( .gnd(gnd), .vdd(vdd), .A(regs_13__20_), .Y(_1843_) );
NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(wdata[20]), .B(_1803__bF_buf7), .Y(_1844_) );
OAI21X1 OAI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_1843_), .B(_1803__bF_buf6), .C(_1844_), .Y(_140_) );
INVX2 INVX2_182 ( .gnd(gnd), .vdd(vdd), .A(regs_13__21_), .Y(_1845_) );
NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(wdata[21]), .B(_1803__bF_buf5), .Y(_1846_) );
OAI21X1 OAI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_1845_), .B(_1803__bF_buf4), .C(_1846_), .Y(_141_) );
INVX2 INVX2_183 ( .gnd(gnd), .vdd(vdd), .A(regs_13__22_), .Y(_1847_) );
NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(wdata[22]), .B(_1803__bF_buf3), .Y(_1848_) );
OAI21X1 OAI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_1847_), .B(_1803__bF_buf2), .C(_1848_), .Y(_142_) );
INVX2 INVX2_184 ( .gnd(gnd), .vdd(vdd), .A(regs_13__23_), .Y(_1849_) );
NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(wdata[23]), .B(_1803__bF_buf1), .Y(_1850_) );
OAI21X1 OAI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_1849_), .B(_1803__bF_buf0), .C(_1850_), .Y(_143_) );
INVX2 INVX2_185 ( .gnd(gnd), .vdd(vdd), .A(regs_13__24_), .Y(_1851_) );
NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(wdata[24]), .B(_1803__bF_buf7), .Y(_1852_) );
OAI21X1 OAI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_1851_), .B(_1803__bF_buf6), .C(_1852_), .Y(_144_) );
INVX2 INVX2_186 ( .gnd(gnd), .vdd(vdd), .A(regs_13__25_), .Y(_1853_) );
NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(wdata[25]), .B(_1803__bF_buf5), .Y(_1854_) );
OAI21X1 OAI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_1853_), .B(_1803__bF_buf4), .C(_1854_), .Y(_145_) );
INVX2 INVX2_187 ( .gnd(gnd), .vdd(vdd), .A(regs_13__26_), .Y(_1855_) );
NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(wdata[26]), .B(_1803__bF_buf3), .Y(_1856_) );
OAI21X1 OAI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_1855_), .B(_1803__bF_buf2), .C(_1856_), .Y(_146_) );
INVX2 INVX2_188 ( .gnd(gnd), .vdd(vdd), .A(regs_13__27_), .Y(_1857_) );
NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(wdata[27]), .B(_1803__bF_buf1), .Y(_1858_) );
OAI21X1 OAI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_1857_), .B(_1803__bF_buf0), .C(_1858_), .Y(_147_) );
INVX2 INVX2_189 ( .gnd(gnd), .vdd(vdd), .A(regs_13__28_), .Y(_1859_) );
NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(wdata[28]), .B(_1803__bF_buf7), .Y(_1860_) );
OAI21X1 OAI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_1859_), .B(_1803__bF_buf6), .C(_1860_), .Y(_148_) );
INVX2 INVX2_190 ( .gnd(gnd), .vdd(vdd), .A(regs_13__29_), .Y(_1861_) );
NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(wdata[29]), .B(_1803__bF_buf5), .Y(_1862_) );
OAI21X1 OAI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_1861_), .B(_1803__bF_buf4), .C(_1862_), .Y(_149_) );
INVX2 INVX2_191 ( .gnd(gnd), .vdd(vdd), .A(regs_13__30_), .Y(_1863_) );
NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(wdata[30]), .B(_1803__bF_buf3), .Y(_1864_) );
OAI21X1 OAI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_1863_), .B(_1803__bF_buf2), .C(_1864_), .Y(_151_) );
INVX2 INVX2_192 ( .gnd(gnd), .vdd(vdd), .A(regs_13__31_), .Y(_1865_) );
NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(wdata[31]), .B(_1803__bF_buf1), .Y(_1866_) );
OAI21X1 OAI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_1865_), .B(_1803__bF_buf0), .C(_1866_), .Y(_152_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf2), .B(_1104__bF_buf10), .Y(_1867_) );
OAI21X1 OAI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf1), .B(_1104__bF_buf9), .C(regs_12__0_), .Y(_1868_) );
OAI21X1 OAI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf4), .B(_992__bF_buf2), .C(_1868_), .Y(_96_) );
OAI21X1 OAI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf0), .B(_1104__bF_buf8), .C(regs_12__1_), .Y(_1869_) );
OAI21X1 OAI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf3), .B(_1003__bF_buf2), .C(_1869_), .Y(_107_) );
OAI21X1 OAI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf5), .B(_1104__bF_buf7), .C(regs_12__2_), .Y(_1870_) );
OAI21X1 OAI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf2), .B(_1005__bF_buf2), .C(_1870_), .Y(_118_) );
OAI21X1 OAI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf4), .B(_1104__bF_buf6), .C(regs_12__3_), .Y(_1871_) );
OAI21X1 OAI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf1), .B(_1007__bF_buf2), .C(_1871_), .Y(_121_) );
OAI21X1 OAI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf3), .B(_1104__bF_buf5), .C(regs_12__4_), .Y(_1872_) );
OAI21X1 OAI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf0), .B(_1009__bF_buf1), .C(_1872_), .Y(_122_) );
OAI21X1 OAI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf2), .B(_1104__bF_buf4), .C(regs_12__5_), .Y(_1873_) );
OAI21X1 OAI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf4), .B(_1011__bF_buf1), .C(_1873_), .Y(_123_) );
OAI21X1 OAI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf1), .B(_1104__bF_buf3), .C(regs_12__6_), .Y(_1874_) );
OAI21X1 OAI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf3), .B(_1013__bF_buf1), .C(_1874_), .Y(_124_) );
OAI21X1 OAI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf0), .B(_1104__bF_buf2), .C(regs_12__7_), .Y(_1875_) );
OAI21X1 OAI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf2), .B(_1015__bF_buf1), .C(_1875_), .Y(_125_) );
OAI21X1 OAI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf5), .B(_1104__bF_buf1), .C(regs_12__8_), .Y(_1876_) );
OAI21X1 OAI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf1), .B(_1017__bF_buf1), .C(_1876_), .Y(_126_) );
OAI21X1 OAI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf4), .B(_1104__bF_buf0), .C(regs_12__9_), .Y(_1877_) );
OAI21X1 OAI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf0), .B(_1019__bF_buf1), .C(_1877_), .Y(_127_) );
OAI21X1 OAI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf3), .B(_1104__bF_buf14), .C(regs_12__10_), .Y(_1878_) );
OAI21X1 OAI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf4), .B(_1021__bF_buf1), .C(_1878_), .Y(_97_) );
OAI21X1 OAI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf2), .B(_1104__bF_buf13), .C(regs_12__11_), .Y(_1879_) );
OAI21X1 OAI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf3), .B(_1023__bF_buf1), .C(_1879_), .Y(_98_) );
OAI21X1 OAI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf1), .B(_1104__bF_buf12), .C(regs_12__12_), .Y(_1880_) );
OAI21X1 OAI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf2), .B(_1025__bF_buf1), .C(_1880_), .Y(_99_) );
OAI21X1 OAI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf0), .B(_1104__bF_buf11), .C(regs_12__13_), .Y(_1881_) );
OAI21X1 OAI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf1), .B(_1027__bF_buf1), .C(_1881_), .Y(_100_) );
OAI21X1 OAI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf5), .B(_1104__bF_buf10), .C(regs_12__14_), .Y(_1882_) );
OAI21X1 OAI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf0), .B(_1029__bF_buf1), .C(_1882_), .Y(_101_) );
OAI21X1 OAI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf4), .B(_1104__bF_buf9), .C(regs_12__15_), .Y(_1883_) );
OAI21X1 OAI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf4), .B(_1031__bF_buf1), .C(_1883_), .Y(_102_) );
OAI21X1 OAI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf3), .B(_1104__bF_buf8), .C(regs_12__16_), .Y(_1884_) );
OAI21X1 OAI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf3), .B(_1033__bF_buf1), .C(_1884_), .Y(_103_) );
OAI21X1 OAI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf2), .B(_1104__bF_buf7), .C(regs_12__17_), .Y(_1885_) );
OAI21X1 OAI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf2), .B(_1035__bF_buf1), .C(_1885_), .Y(_104_) );
OAI21X1 OAI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf1), .B(_1104__bF_buf6), .C(regs_12__18_), .Y(_1886_) );
OAI21X1 OAI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf1), .B(_1037__bF_buf1), .C(_1886_), .Y(_105_) );
OAI21X1 OAI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf0), .B(_1104__bF_buf5), .C(regs_12__19_), .Y(_1887_) );
OAI21X1 OAI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf0), .B(_1039__bF_buf1), .C(_1887_), .Y(_106_) );
OAI21X1 OAI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf5), .B(_1104__bF_buf4), .C(regs_12__20_), .Y(_1888_) );
OAI21X1 OAI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf4), .B(_1041__bF_buf1), .C(_1888_), .Y(_108_) );
OAI21X1 OAI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf4), .B(_1104__bF_buf3), .C(regs_12__21_), .Y(_1889_) );
OAI21X1 OAI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf3), .B(_1043__bF_buf1), .C(_1889_), .Y(_109_) );
OAI21X1 OAI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf3), .B(_1104__bF_buf2), .C(regs_12__22_), .Y(_1890_) );
OAI21X1 OAI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf2), .B(_1045__bF_buf1), .C(_1890_), .Y(_110_) );
OAI21X1 OAI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf2), .B(_1104__bF_buf1), .C(regs_12__23_), .Y(_1891_) );
OAI21X1 OAI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf1), .B(_1047__bF_buf1), .C(_1891_), .Y(_111_) );
OAI21X1 OAI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf1), .B(_1104__bF_buf0), .C(regs_12__24_), .Y(_1892_) );
OAI21X1 OAI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf0), .B(_1049__bF_buf1), .C(_1892_), .Y(_112_) );
OAI21X1 OAI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf0), .B(_1104__bF_buf14), .C(regs_12__25_), .Y(_1893_) );
OAI21X1 OAI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf4), .B(_1051__bF_buf1), .C(_1893_), .Y(_113_) );
OAI21X1 OAI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf5), .B(_1104__bF_buf13), .C(regs_12__26_), .Y(_1894_) );
OAI21X1 OAI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf3), .B(_1053__bF_buf1), .C(_1894_), .Y(_114_) );
OAI21X1 OAI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf4), .B(_1104__bF_buf12), .C(regs_12__27_), .Y(_1895_) );
OAI21X1 OAI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf2), .B(_1055__bF_buf1), .C(_1895_), .Y(_115_) );
OAI21X1 OAI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf3), .B(_1104__bF_buf11), .C(regs_12__28_), .Y(_1896_) );
OAI21X1 OAI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf1), .B(_1057__bF_buf1), .C(_1896_), .Y(_116_) );
OAI21X1 OAI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf2), .B(_1104__bF_buf10), .C(regs_12__29_), .Y(_1897_) );
OAI21X1 OAI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf0), .B(_1059__bF_buf1), .C(_1897_), .Y(_117_) );
OAI21X1 OAI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf1), .B(_1104__bF_buf9), .C(regs_12__30_), .Y(_1898_) );
OAI21X1 OAI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf4), .B(_1061__bF_buf1), .C(_1898_), .Y(_119_) );
OAI21X1 OAI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(_1704__bF_buf0), .B(_1104__bF_buf8), .C(regs_12__31_), .Y(_1899_) );
OAI21X1 OAI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(_1867__bF_buf3), .B(_1063__bF_buf1), .C(_1899_), .Y(_120_) );
INVX2 INVX2_193 ( .gnd(gnd), .vdd(vdd), .A(regs_11__0_), .Y(_1900_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_1703_), .B(_1139_), .Y(_1901_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1142__bF_buf2), .B(_1901__bF_buf5), .Y(_1902_) );
NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(wdata[0]), .B(_1902__bF_buf7), .Y(_1903_) );
OAI21X1 OAI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(_1900_), .B(_1902__bF_buf6), .C(_1903_), .Y(_64_) );
INVX2 INVX2_194 ( .gnd(gnd), .vdd(vdd), .A(regs_11__1_), .Y(_1904_) );
NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(wdata[1]), .B(_1902__bF_buf5), .Y(_1905_) );
OAI21X1 OAI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(_1904_), .B(_1902__bF_buf4), .C(_1905_), .Y(_75_) );
INVX2 INVX2_195 ( .gnd(gnd), .vdd(vdd), .A(regs_11__2_), .Y(_1906_) );
NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(wdata[2]), .B(_1902__bF_buf3), .Y(_1907_) );
OAI21X1 OAI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_1906_), .B(_1902__bF_buf2), .C(_1907_), .Y(_86_) );
INVX2 INVX2_196 ( .gnd(gnd), .vdd(vdd), .A(regs_11__3_), .Y(_1908_) );
NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(wdata[3]), .B(_1902__bF_buf1), .Y(_1909_) );
OAI21X1 OAI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_1908_), .B(_1902__bF_buf0), .C(_1909_), .Y(_89_) );
INVX2 INVX2_197 ( .gnd(gnd), .vdd(vdd), .A(regs_11__4_), .Y(_1910_) );
NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(wdata[4]), .B(_1902__bF_buf7), .Y(_1911_) );
OAI21X1 OAI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(_1910_), .B(_1902__bF_buf6), .C(_1911_), .Y(_90_) );
INVX2 INVX2_198 ( .gnd(gnd), .vdd(vdd), .A(regs_11__5_), .Y(_1912_) );
NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(wdata[5]), .B(_1902__bF_buf5), .Y(_1913_) );
OAI21X1 OAI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(_1912_), .B(_1902__bF_buf4), .C(_1913_), .Y(_91_) );
INVX2 INVX2_199 ( .gnd(gnd), .vdd(vdd), .A(regs_11__6_), .Y(_1914_) );
NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(wdata[6]), .B(_1902__bF_buf3), .Y(_1915_) );
OAI21X1 OAI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_1914_), .B(_1902__bF_buf2), .C(_1915_), .Y(_92_) );
INVX2 INVX2_200 ( .gnd(gnd), .vdd(vdd), .A(regs_11__7_), .Y(_1916_) );
NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(wdata[7]), .B(_1902__bF_buf1), .Y(_1917_) );
OAI21X1 OAI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(_1916_), .B(_1902__bF_buf0), .C(_1917_), .Y(_93_) );
INVX2 INVX2_201 ( .gnd(gnd), .vdd(vdd), .A(regs_11__8_), .Y(_1918_) );
NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(wdata[8]), .B(_1902__bF_buf7), .Y(_1919_) );
OAI21X1 OAI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_1918_), .B(_1902__bF_buf6), .C(_1919_), .Y(_94_) );
INVX2 INVX2_202 ( .gnd(gnd), .vdd(vdd), .A(regs_11__9_), .Y(_1920_) );
NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(wdata[9]), .B(_1902__bF_buf5), .Y(_1921_) );
OAI21X1 OAI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_1920_), .B(_1902__bF_buf4), .C(_1921_), .Y(_95_) );
INVX2 INVX2_203 ( .gnd(gnd), .vdd(vdd), .A(regs_11__10_), .Y(_1922_) );
NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(wdata[10]), .B(_1902__bF_buf3), .Y(_1923_) );
OAI21X1 OAI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_1922_), .B(_1902__bF_buf2), .C(_1923_), .Y(_65_) );
INVX2 INVX2_204 ( .gnd(gnd), .vdd(vdd), .A(regs_11__11_), .Y(_1924_) );
NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(wdata[11]), .B(_1902__bF_buf1), .Y(_1925_) );
OAI21X1 OAI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_1924_), .B(_1902__bF_buf0), .C(_1925_), .Y(_66_) );
INVX2 INVX2_205 ( .gnd(gnd), .vdd(vdd), .A(regs_11__12_), .Y(_1926_) );
NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(wdata[12]), .B(_1902__bF_buf7), .Y(_1927_) );
OAI21X1 OAI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_1926_), .B(_1902__bF_buf6), .C(_1927_), .Y(_67_) );
INVX2 INVX2_206 ( .gnd(gnd), .vdd(vdd), .A(regs_11__13_), .Y(_1928_) );
NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(wdata[13]), .B(_1902__bF_buf5), .Y(_1929_) );
OAI21X1 OAI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_1928_), .B(_1902__bF_buf4), .C(_1929_), .Y(_68_) );
INVX2 INVX2_207 ( .gnd(gnd), .vdd(vdd), .A(regs_11__14_), .Y(_1930_) );
NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(wdata[14]), .B(_1902__bF_buf3), .Y(_1931_) );
OAI21X1 OAI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_1930_), .B(_1902__bF_buf2), .C(_1931_), .Y(_69_) );
INVX2 INVX2_208 ( .gnd(gnd), .vdd(vdd), .A(regs_11__15_), .Y(_1932_) );
NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(wdata[15]), .B(_1902__bF_buf1), .Y(_1933_) );
OAI21X1 OAI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_1932_), .B(_1902__bF_buf0), .C(_1933_), .Y(_70_) );
INVX2 INVX2_209 ( .gnd(gnd), .vdd(vdd), .A(regs_11__16_), .Y(_1934_) );
NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(wdata[16]), .B(_1902__bF_buf7), .Y(_1935_) );
OAI21X1 OAI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_1934_), .B(_1902__bF_buf6), .C(_1935_), .Y(_71_) );
INVX2 INVX2_210 ( .gnd(gnd), .vdd(vdd), .A(regs_11__17_), .Y(_1936_) );
NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(wdata[17]), .B(_1902__bF_buf5), .Y(_1937_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_5511__0_), .Y(rdata1[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_5511__1_), .Y(rdata1[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_5511__2_), .Y(rdata1[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_5511__3_), .Y(rdata1[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_5511__4_), .Y(rdata1[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_5511__5_), .Y(rdata1[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_5511__6_), .Y(rdata1[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_5511__7_), .Y(rdata1[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_5511__8_), .Y(rdata1[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_5511__9_), .Y(rdata1[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_5511__10_), .Y(rdata1[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_5511__11_), .Y(rdata1[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_5511__12_), .Y(rdata1[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_5511__13_), .Y(rdata1[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_5511__14_), .Y(rdata1[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_5511__15_), .Y(rdata1[15]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_5511__16_), .Y(rdata1[16]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_5511__17_), .Y(rdata1[17]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_5511__18_), .Y(rdata1[18]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_5511__19_), .Y(rdata1[19]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_5511__20_), .Y(rdata1[20]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_5511__21_), .Y(rdata1[21]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_5511__22_), .Y(rdata1[22]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_5511__23_), .Y(rdata1[23]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_5511__24_), .Y(rdata1[24]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_5511__25_), .Y(rdata1[25]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_5511__26_), .Y(rdata1[26]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_5511__27_), .Y(rdata1[27]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_5511__28_), .Y(rdata1[28]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_5511__29_), .Y(rdata1[29]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_5511__30_), .Y(rdata1[30]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_5511__31_), .Y(rdata1[31]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_5512__0_), .Y(rdata2[0]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_5512__1_), .Y(rdata2[1]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_5512__2_), .Y(rdata2[2]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_5512__3_), .Y(rdata2[3]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_5512__4_), .Y(rdata2[4]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_5512__5_), .Y(rdata2[5]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_5512__6_), .Y(rdata2[6]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_5512__7_), .Y(rdata2[7]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_5512__8_), .Y(rdata2[8]) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_5512__9_), .Y(rdata2[9]) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_5512__10_), .Y(rdata2[10]) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_5512__11_), .Y(rdata2[11]) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_5512__12_), .Y(rdata2[12]) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_5512__13_), .Y(rdata2[13]) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_5512__14_), .Y(rdata2[14]) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(_5512__15_), .Y(rdata2[15]) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(_5512__16_), .Y(rdata2[16]) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(_5512__17_), .Y(rdata2[17]) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(_5512__18_), .Y(rdata2[18]) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(_5512__19_), .Y(rdata2[19]) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(_5512__20_), .Y(rdata2[20]) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(_5512__21_), .Y(rdata2[21]) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(_5512__22_), .Y(rdata2[22]) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(_5512__23_), .Y(rdata2[23]) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(_5512__24_), .Y(rdata2[24]) );
BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(_5512__25_), .Y(rdata2[25]) );
BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(_5512__26_), .Y(rdata2[26]) );
BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(_5512__27_), .Y(rdata2[27]) );
BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(_5512__28_), .Y(rdata2[28]) );
BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(_5512__29_), .Y(rdata2[29]) );
BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(_5512__30_), .Y(rdata2[30]) );
BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(_5512__31_), .Y(rdata2[31]) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_352_), .Q(regs_1__0_) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_363_), .Q(regs_1__1_) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_374_), .Q(regs_1__2_) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_377_), .Q(regs_1__3_) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_378_), .Q(regs_1__4_) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_379_), .Q(regs_1__5_) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_380_), .Q(regs_1__6_) );
DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_381_), .Q(regs_1__7_) );
DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_382_), .Q(regs_1__8_) );
DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_383_), .Q(regs_1__9_) );
DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_353_), .Q(regs_1__10_) );
DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_354_), .Q(regs_1__11_) );
DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_355_), .Q(regs_1__12_) );
DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_356_), .Q(regs_1__13_) );
DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_357_), .Q(regs_1__14_) );
DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_358_), .Q(regs_1__15_) );
DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_359_), .Q(regs_1__16_) );
DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_360_), .Q(regs_1__17_) );
DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_361_), .Q(regs_1__18_) );
DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_362_), .Q(regs_1__19_) );
DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_364_), .Q(regs_1__20_) );
DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_365_), .Q(regs_1__21_) );
DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_366_), .Q(regs_1__22_) );
DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_367_), .Q(regs_1__23_) );
DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_368_), .Q(regs_1__24_) );
DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_369_), .Q(regs_1__25_) );
DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_370_), .Q(regs_1__26_) );
DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_371_), .Q(regs_1__27_) );
DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_372_), .Q(regs_1__28_) );
DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_373_), .Q(regs_1__29_) );
DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_375_), .Q(regs_1__30_) );
DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_376_), .Q(regs_1__31_) );
DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_0_), .Q(regs_0__0_) );
DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_11_), .Q(regs_0__1_) );
DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_22_), .Q(regs_0__2_) );
DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_25_), .Q(regs_0__3_) );
DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_26_), .Q(regs_0__4_) );
DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_27_), .Q(regs_0__5_) );
DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_28_), .Q(regs_0__6_) );
DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_29_), .Q(regs_0__7_) );
DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_30_), .Q(regs_0__8_) );
DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_31_), .Q(regs_0__9_) );
DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_1_), .Q(regs_0__10_) );
DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_2_), .Q(regs_0__11_) );
DFFPOSX1 DFFPOSX1_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_3_), .Q(regs_0__12_) );
DFFPOSX1 DFFPOSX1_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_4_), .Q(regs_0__13_) );
DFFPOSX1 DFFPOSX1_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_5_), .Q(regs_0__14_) );
DFFPOSX1 DFFPOSX1_48 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_6_), .Q(regs_0__15_) );
DFFPOSX1 DFFPOSX1_49 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_7_), .Q(regs_0__16_) );
DFFPOSX1 DFFPOSX1_50 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_8_), .Q(regs_0__17_) );
DFFPOSX1 DFFPOSX1_51 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_9_), .Q(regs_0__18_) );
DFFPOSX1 DFFPOSX1_52 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_10_), .Q(regs_0__19_) );
DFFPOSX1 DFFPOSX1_53 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_12_), .Q(regs_0__20_) );
DFFPOSX1 DFFPOSX1_54 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_13_), .Q(regs_0__21_) );
DFFPOSX1 DFFPOSX1_55 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_14_), .Q(regs_0__22_) );
DFFPOSX1 DFFPOSX1_56 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_15_), .Q(regs_0__23_) );
DFFPOSX1 DFFPOSX1_57 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_16_), .Q(regs_0__24_) );
DFFPOSX1 DFFPOSX1_58 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_17_), .Q(regs_0__25_) );
DFFPOSX1 DFFPOSX1_59 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_18_), .Q(regs_0__26_) );
DFFPOSX1 DFFPOSX1_60 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_19_), .Q(regs_0__27_) );
DFFPOSX1 DFFPOSX1_61 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_20_), .Q(regs_0__28_) );
DFFPOSX1 DFFPOSX1_62 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_21_), .Q(regs_0__29_) );
DFFPOSX1 DFFPOSX1_63 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_23_), .Q(regs_0__30_) );
DFFPOSX1 DFFPOSX1_64 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_24_), .Q(regs_0__31_) );
DFFPOSX1 DFFPOSX1_65 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_640_), .Q(regs_28__0_) );
DFFPOSX1 DFFPOSX1_66 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_651_), .Q(regs_28__1_) );
DFFPOSX1 DFFPOSX1_67 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_662_), .Q(regs_28__2_) );
DFFPOSX1 DFFPOSX1_68 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_665_), .Q(regs_28__3_) );
DFFPOSX1 DFFPOSX1_69 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_666_), .Q(regs_28__4_) );
DFFPOSX1 DFFPOSX1_70 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_667_), .Q(regs_28__5_) );
DFFPOSX1 DFFPOSX1_71 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_668_), .Q(regs_28__6_) );
DFFPOSX1 DFFPOSX1_72 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_669_), .Q(regs_28__7_) );
DFFPOSX1 DFFPOSX1_73 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_670_), .Q(regs_28__8_) );
DFFPOSX1 DFFPOSX1_74 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_671_), .Q(regs_28__9_) );
DFFPOSX1 DFFPOSX1_75 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_641_), .Q(regs_28__10_) );
DFFPOSX1 DFFPOSX1_76 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_642_), .Q(regs_28__11_) );
DFFPOSX1 DFFPOSX1_77 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_643_), .Q(regs_28__12_) );
DFFPOSX1 DFFPOSX1_78 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_644_), .Q(regs_28__13_) );
DFFPOSX1 DFFPOSX1_79 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_645_), .Q(regs_28__14_) );
DFFPOSX1 DFFPOSX1_80 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_646_), .Q(regs_28__15_) );
DFFPOSX1 DFFPOSX1_81 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_647_), .Q(regs_28__16_) );
DFFPOSX1 DFFPOSX1_82 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_648_), .Q(regs_28__17_) );
DFFPOSX1 DFFPOSX1_83 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_649_), .Q(regs_28__18_) );
DFFPOSX1 DFFPOSX1_84 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_650_), .Q(regs_28__19_) );
DFFPOSX1 DFFPOSX1_85 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_652_), .Q(regs_28__20_) );
DFFPOSX1 DFFPOSX1_86 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_653_), .Q(regs_28__21_) );
DFFPOSX1 DFFPOSX1_87 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_654_), .Q(regs_28__22_) );
DFFPOSX1 DFFPOSX1_88 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_655_), .Q(regs_28__23_) );
DFFPOSX1 DFFPOSX1_89 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_656_), .Q(regs_28__24_) );
DFFPOSX1 DFFPOSX1_90 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_657_), .Q(regs_28__25_) );
DFFPOSX1 DFFPOSX1_91 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_658_), .Q(regs_28__26_) );
DFFPOSX1 DFFPOSX1_92 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_659_), .Q(regs_28__27_) );
DFFPOSX1 DFFPOSX1_93 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_660_), .Q(regs_28__28_) );
DFFPOSX1 DFFPOSX1_94 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_661_), .Q(regs_28__29_) );
DFFPOSX1 DFFPOSX1_95 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_663_), .Q(regs_28__30_) );
DFFPOSX1 DFFPOSX1_96 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_664_), .Q(regs_28__31_) );
DFFPOSX1 DFFPOSX1_97 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_736_), .Q(regs_30__0_) );
DFFPOSX1 DFFPOSX1_98 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_747_), .Q(regs_30__1_) );
DFFPOSX1 DFFPOSX1_99 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_758_), .Q(regs_30__2_) );
DFFPOSX1 DFFPOSX1_100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_761_), .Q(regs_30__3_) );
DFFPOSX1 DFFPOSX1_101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_762_), .Q(regs_30__4_) );
DFFPOSX1 DFFPOSX1_102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_763_), .Q(regs_30__5_) );
DFFPOSX1 DFFPOSX1_103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_764_), .Q(regs_30__6_) );
DFFPOSX1 DFFPOSX1_104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_765_), .Q(regs_30__7_) );
DFFPOSX1 DFFPOSX1_105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_766_), .Q(regs_30__8_) );
DFFPOSX1 DFFPOSX1_106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_767_), .Q(regs_30__9_) );
DFFPOSX1 DFFPOSX1_107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_737_), .Q(regs_30__10_) );
DFFPOSX1 DFFPOSX1_108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_738_), .Q(regs_30__11_) );
DFFPOSX1 DFFPOSX1_109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_739_), .Q(regs_30__12_) );
DFFPOSX1 DFFPOSX1_110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_740_), .Q(regs_30__13_) );
DFFPOSX1 DFFPOSX1_111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_741_), .Q(regs_30__14_) );
DFFPOSX1 DFFPOSX1_112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_742_), .Q(regs_30__15_) );
DFFPOSX1 DFFPOSX1_113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_743_), .Q(regs_30__16_) );
DFFPOSX1 DFFPOSX1_114 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_744_), .Q(regs_30__17_) );
DFFPOSX1 DFFPOSX1_115 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_745_), .Q(regs_30__18_) );
DFFPOSX1 DFFPOSX1_116 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_746_), .Q(regs_30__19_) );
DFFPOSX1 DFFPOSX1_117 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_748_), .Q(regs_30__20_) );
DFFPOSX1 DFFPOSX1_118 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_749_), .Q(regs_30__21_) );
DFFPOSX1 DFFPOSX1_119 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_750_), .Q(regs_30__22_) );
DFFPOSX1 DFFPOSX1_120 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_751_), .Q(regs_30__23_) );
DFFPOSX1 DFFPOSX1_121 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_752_), .Q(regs_30__24_) );
DFFPOSX1 DFFPOSX1_122 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_753_), .Q(regs_30__25_) );
DFFPOSX1 DFFPOSX1_123 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_754_), .Q(regs_30__26_) );
DFFPOSX1 DFFPOSX1_124 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_755_), .Q(regs_30__27_) );
DFFPOSX1 DFFPOSX1_125 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_756_), .Q(regs_30__28_) );
DFFPOSX1 DFFPOSX1_126 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_757_), .Q(regs_30__29_) );
DFFPOSX1 DFFPOSX1_127 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_759_), .Q(regs_30__30_) );
DFFPOSX1 DFFPOSX1_128 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_760_), .Q(regs_30__31_) );
DFFPOSX1 DFFPOSX1_129 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_672_), .Q(regs_29__0_) );
DFFPOSX1 DFFPOSX1_130 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_683_), .Q(regs_29__1_) );
DFFPOSX1 DFFPOSX1_131 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_694_), .Q(regs_29__2_) );
DFFPOSX1 DFFPOSX1_132 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_697_), .Q(regs_29__3_) );
DFFPOSX1 DFFPOSX1_133 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_698_), .Q(regs_29__4_) );
DFFPOSX1 DFFPOSX1_134 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_699_), .Q(regs_29__5_) );
DFFPOSX1 DFFPOSX1_135 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_700_), .Q(regs_29__6_) );
DFFPOSX1 DFFPOSX1_136 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_701_), .Q(regs_29__7_) );
DFFPOSX1 DFFPOSX1_137 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_702_), .Q(regs_29__8_) );
DFFPOSX1 DFFPOSX1_138 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_703_), .Q(regs_29__9_) );
DFFPOSX1 DFFPOSX1_139 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_673_), .Q(regs_29__10_) );
DFFPOSX1 DFFPOSX1_140 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_674_), .Q(regs_29__11_) );
DFFPOSX1 DFFPOSX1_141 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_675_), .Q(regs_29__12_) );
DFFPOSX1 DFFPOSX1_142 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_676_), .Q(regs_29__13_) );
DFFPOSX1 DFFPOSX1_143 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_677_), .Q(regs_29__14_) );
DFFPOSX1 DFFPOSX1_144 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_678_), .Q(regs_29__15_) );
DFFPOSX1 DFFPOSX1_145 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_679_), .Q(regs_29__16_) );
DFFPOSX1 DFFPOSX1_146 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_680_), .Q(regs_29__17_) );
DFFPOSX1 DFFPOSX1_147 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_681_), .Q(regs_29__18_) );
DFFPOSX1 DFFPOSX1_148 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_682_), .Q(regs_29__19_) );
DFFPOSX1 DFFPOSX1_149 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_684_), .Q(regs_29__20_) );
DFFPOSX1 DFFPOSX1_150 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_685_), .Q(regs_29__21_) );
DFFPOSX1 DFFPOSX1_151 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_686_), .Q(regs_29__22_) );
DFFPOSX1 DFFPOSX1_152 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_687_), .Q(regs_29__23_) );
DFFPOSX1 DFFPOSX1_153 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_688_), .Q(regs_29__24_) );
DFFPOSX1 DFFPOSX1_154 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_689_), .Q(regs_29__25_) );
DFFPOSX1 DFFPOSX1_155 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_690_), .Q(regs_29__26_) );
DFFPOSX1 DFFPOSX1_156 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_691_), .Q(regs_29__27_) );
DFFPOSX1 DFFPOSX1_157 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_692_), .Q(regs_29__28_) );
DFFPOSX1 DFFPOSX1_158 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_693_), .Q(regs_29__29_) );
DFFPOSX1 DFFPOSX1_159 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_695_), .Q(regs_29__30_) );
DFFPOSX1 DFFPOSX1_160 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_696_), .Q(regs_29__31_) );
DFFPOSX1 DFFPOSX1_161 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_608_), .Q(regs_27__0_) );
DFFPOSX1 DFFPOSX1_162 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_619_), .Q(regs_27__1_) );
DFFPOSX1 DFFPOSX1_163 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_630_), .Q(regs_27__2_) );
DFFPOSX1 DFFPOSX1_164 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_633_), .Q(regs_27__3_) );
DFFPOSX1 DFFPOSX1_165 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_634_), .Q(regs_27__4_) );
DFFPOSX1 DFFPOSX1_166 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_635_), .Q(regs_27__5_) );
DFFPOSX1 DFFPOSX1_167 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_636_), .Q(regs_27__6_) );
DFFPOSX1 DFFPOSX1_168 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_637_), .Q(regs_27__7_) );
DFFPOSX1 DFFPOSX1_169 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_638_), .Q(regs_27__8_) );
DFFPOSX1 DFFPOSX1_170 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_639_), .Q(regs_27__9_) );
DFFPOSX1 DFFPOSX1_171 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_609_), .Q(regs_27__10_) );
DFFPOSX1 DFFPOSX1_172 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_610_), .Q(regs_27__11_) );
DFFPOSX1 DFFPOSX1_173 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_611_), .Q(regs_27__12_) );
DFFPOSX1 DFFPOSX1_174 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_612_), .Q(regs_27__13_) );
DFFPOSX1 DFFPOSX1_175 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_613_), .Q(regs_27__14_) );
DFFPOSX1 DFFPOSX1_176 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_614_), .Q(regs_27__15_) );
DFFPOSX1 DFFPOSX1_177 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_615_), .Q(regs_27__16_) );
DFFPOSX1 DFFPOSX1_178 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_616_), .Q(regs_27__17_) );
DFFPOSX1 DFFPOSX1_179 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_617_), .Q(regs_27__18_) );
DFFPOSX1 DFFPOSX1_180 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_618_), .Q(regs_27__19_) );
DFFPOSX1 DFFPOSX1_181 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_620_), .Q(regs_27__20_) );
DFFPOSX1 DFFPOSX1_182 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_621_), .Q(regs_27__21_) );
DFFPOSX1 DFFPOSX1_183 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_622_), .Q(regs_27__22_) );
DFFPOSX1 DFFPOSX1_184 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_623_), .Q(regs_27__23_) );
DFFPOSX1 DFFPOSX1_185 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_624_), .Q(regs_27__24_) );
DFFPOSX1 DFFPOSX1_186 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_625_), .Q(regs_27__25_) );
DFFPOSX1 DFFPOSX1_187 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_626_), .Q(regs_27__26_) );
DFFPOSX1 DFFPOSX1_188 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_627_), .Q(regs_27__27_) );
DFFPOSX1 DFFPOSX1_189 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_628_), .Q(regs_27__28_) );
DFFPOSX1 DFFPOSX1_190 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_629_), .Q(regs_27__29_) );
DFFPOSX1 DFFPOSX1_191 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_631_), .Q(regs_27__30_) );
DFFPOSX1 DFFPOSX1_192 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_632_), .Q(regs_27__31_) );
DFFPOSX1 DFFPOSX1_193 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_576_), .Q(regs_26__0_) );
DFFPOSX1 DFFPOSX1_194 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_587_), .Q(regs_26__1_) );
DFFPOSX1 DFFPOSX1_195 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_598_), .Q(regs_26__2_) );
DFFPOSX1 DFFPOSX1_196 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_601_), .Q(regs_26__3_) );
DFFPOSX1 DFFPOSX1_197 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_602_), .Q(regs_26__4_) );
DFFPOSX1 DFFPOSX1_198 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_603_), .Q(regs_26__5_) );
DFFPOSX1 DFFPOSX1_199 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_604_), .Q(regs_26__6_) );
DFFPOSX1 DFFPOSX1_200 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_605_), .Q(regs_26__7_) );
DFFPOSX1 DFFPOSX1_201 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_606_), .Q(regs_26__8_) );
DFFPOSX1 DFFPOSX1_202 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_607_), .Q(regs_26__9_) );
DFFPOSX1 DFFPOSX1_203 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_577_), .Q(regs_26__10_) );
DFFPOSX1 DFFPOSX1_204 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_578_), .Q(regs_26__11_) );
DFFPOSX1 DFFPOSX1_205 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_579_), .Q(regs_26__12_) );
DFFPOSX1 DFFPOSX1_206 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_580_), .Q(regs_26__13_) );
DFFPOSX1 DFFPOSX1_207 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_581_), .Q(regs_26__14_) );
DFFPOSX1 DFFPOSX1_208 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_582_), .Q(regs_26__15_) );
DFFPOSX1 DFFPOSX1_209 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_583_), .Q(regs_26__16_) );
DFFPOSX1 DFFPOSX1_210 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_584_), .Q(regs_26__17_) );
DFFPOSX1 DFFPOSX1_211 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_585_), .Q(regs_26__18_) );
DFFPOSX1 DFFPOSX1_212 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_586_), .Q(regs_26__19_) );
DFFPOSX1 DFFPOSX1_213 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_588_), .Q(regs_26__20_) );
DFFPOSX1 DFFPOSX1_214 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_589_), .Q(regs_26__21_) );
DFFPOSX1 DFFPOSX1_215 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_590_), .Q(regs_26__22_) );
DFFPOSX1 DFFPOSX1_216 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_591_), .Q(regs_26__23_) );
DFFPOSX1 DFFPOSX1_217 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_592_), .Q(regs_26__24_) );
DFFPOSX1 DFFPOSX1_218 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_593_), .Q(regs_26__25_) );
DFFPOSX1 DFFPOSX1_219 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_594_), .Q(regs_26__26_) );
DFFPOSX1 DFFPOSX1_220 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_595_), .Q(regs_26__27_) );
DFFPOSX1 DFFPOSX1_221 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_596_), .Q(regs_26__28_) );
DFFPOSX1 DFFPOSX1_222 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_597_), .Q(regs_26__29_) );
DFFPOSX1 DFFPOSX1_223 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_599_), .Q(regs_26__30_) );
DFFPOSX1 DFFPOSX1_224 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_600_), .Q(regs_26__31_) );
DFFPOSX1 DFFPOSX1_225 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_544_), .Q(regs_25__0_) );
DFFPOSX1 DFFPOSX1_226 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_555_), .Q(regs_25__1_) );
DFFPOSX1 DFFPOSX1_227 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_566_), .Q(regs_25__2_) );
DFFPOSX1 DFFPOSX1_228 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_569_), .Q(regs_25__3_) );
DFFPOSX1 DFFPOSX1_229 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_570_), .Q(regs_25__4_) );
DFFPOSX1 DFFPOSX1_230 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_571_), .Q(regs_25__5_) );
DFFPOSX1 DFFPOSX1_231 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_572_), .Q(regs_25__6_) );
DFFPOSX1 DFFPOSX1_232 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_573_), .Q(regs_25__7_) );
DFFPOSX1 DFFPOSX1_233 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_574_), .Q(regs_25__8_) );
DFFPOSX1 DFFPOSX1_234 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_575_), .Q(regs_25__9_) );
DFFPOSX1 DFFPOSX1_235 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_545_), .Q(regs_25__10_) );
DFFPOSX1 DFFPOSX1_236 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_546_), .Q(regs_25__11_) );
DFFPOSX1 DFFPOSX1_237 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_547_), .Q(regs_25__12_) );
DFFPOSX1 DFFPOSX1_238 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_548_), .Q(regs_25__13_) );
DFFPOSX1 DFFPOSX1_239 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_549_), .Q(regs_25__14_) );
DFFPOSX1 DFFPOSX1_240 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_550_), .Q(regs_25__15_) );
DFFPOSX1 DFFPOSX1_241 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_551_), .Q(regs_25__16_) );
DFFPOSX1 DFFPOSX1_242 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_552_), .Q(regs_25__17_) );
DFFPOSX1 DFFPOSX1_243 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_553_), .Q(regs_25__18_) );
DFFPOSX1 DFFPOSX1_244 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_554_), .Q(regs_25__19_) );
DFFPOSX1 DFFPOSX1_245 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_556_), .Q(regs_25__20_) );
DFFPOSX1 DFFPOSX1_246 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_557_), .Q(regs_25__21_) );
DFFPOSX1 DFFPOSX1_247 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_558_), .Q(regs_25__22_) );
DFFPOSX1 DFFPOSX1_248 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_559_), .Q(regs_25__23_) );
DFFPOSX1 DFFPOSX1_249 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_560_), .Q(regs_25__24_) );
DFFPOSX1 DFFPOSX1_250 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_561_), .Q(regs_25__25_) );
DFFPOSX1 DFFPOSX1_251 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_562_), .Q(regs_25__26_) );
DFFPOSX1 DFFPOSX1_252 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_563_), .Q(regs_25__27_) );
DFFPOSX1 DFFPOSX1_253 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_564_), .Q(regs_25__28_) );
DFFPOSX1 DFFPOSX1_254 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_565_), .Q(regs_25__29_) );
DFFPOSX1 DFFPOSX1_255 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_567_), .Q(regs_25__30_) );
DFFPOSX1 DFFPOSX1_256 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_568_), .Q(regs_25__31_) );
DFFPOSX1 DFFPOSX1_257 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_512_), .Q(regs_24__0_) );
DFFPOSX1 DFFPOSX1_258 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_523_), .Q(regs_24__1_) );
DFFPOSX1 DFFPOSX1_259 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_534_), .Q(regs_24__2_) );
DFFPOSX1 DFFPOSX1_260 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_537_), .Q(regs_24__3_) );
DFFPOSX1 DFFPOSX1_261 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_538_), .Q(regs_24__4_) );
DFFPOSX1 DFFPOSX1_262 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_539_), .Q(regs_24__5_) );
DFFPOSX1 DFFPOSX1_263 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_540_), .Q(regs_24__6_) );
DFFPOSX1 DFFPOSX1_264 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_541_), .Q(regs_24__7_) );
DFFPOSX1 DFFPOSX1_265 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_542_), .Q(regs_24__8_) );
DFFPOSX1 DFFPOSX1_266 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_543_), .Q(regs_24__9_) );
DFFPOSX1 DFFPOSX1_267 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_513_), .Q(regs_24__10_) );
DFFPOSX1 DFFPOSX1_268 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_514_), .Q(regs_24__11_) );
DFFPOSX1 DFFPOSX1_269 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_515_), .Q(regs_24__12_) );
DFFPOSX1 DFFPOSX1_270 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_516_), .Q(regs_24__13_) );
DFFPOSX1 DFFPOSX1_271 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_517_), .Q(regs_24__14_) );
DFFPOSX1 DFFPOSX1_272 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_518_), .Q(regs_24__15_) );
DFFPOSX1 DFFPOSX1_273 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_519_), .Q(regs_24__16_) );
DFFPOSX1 DFFPOSX1_274 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_520_), .Q(regs_24__17_) );
DFFPOSX1 DFFPOSX1_275 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_521_), .Q(regs_24__18_) );
DFFPOSX1 DFFPOSX1_276 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_522_), .Q(regs_24__19_) );
DFFPOSX1 DFFPOSX1_277 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_524_), .Q(regs_24__20_) );
DFFPOSX1 DFFPOSX1_278 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_525_), .Q(regs_24__21_) );
DFFPOSX1 DFFPOSX1_279 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_526_), .Q(regs_24__22_) );
DFFPOSX1 DFFPOSX1_280 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_527_), .Q(regs_24__23_) );
DFFPOSX1 DFFPOSX1_281 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_528_), .Q(regs_24__24_) );
DFFPOSX1 DFFPOSX1_282 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_529_), .Q(regs_24__25_) );
DFFPOSX1 DFFPOSX1_283 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_530_), .Q(regs_24__26_) );
DFFPOSX1 DFFPOSX1_284 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_531_), .Q(regs_24__27_) );
DFFPOSX1 DFFPOSX1_285 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_532_), .Q(regs_24__28_) );
DFFPOSX1 DFFPOSX1_286 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_533_), .Q(regs_24__29_) );
DFFPOSX1 DFFPOSX1_287 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_535_), .Q(regs_24__30_) );
DFFPOSX1 DFFPOSX1_288 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_536_), .Q(regs_24__31_) );
DFFPOSX1 DFFPOSX1_289 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_480_), .Q(regs_23__0_) );
DFFPOSX1 DFFPOSX1_290 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_491_), .Q(regs_23__1_) );
DFFPOSX1 DFFPOSX1_291 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_502_), .Q(regs_23__2_) );
DFFPOSX1 DFFPOSX1_292 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_505_), .Q(regs_23__3_) );
DFFPOSX1 DFFPOSX1_293 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_506_), .Q(regs_23__4_) );
DFFPOSX1 DFFPOSX1_294 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_507_), .Q(regs_23__5_) );
DFFPOSX1 DFFPOSX1_295 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_508_), .Q(regs_23__6_) );
DFFPOSX1 DFFPOSX1_296 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_509_), .Q(regs_23__7_) );
DFFPOSX1 DFFPOSX1_297 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_510_), .Q(regs_23__8_) );
DFFPOSX1 DFFPOSX1_298 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_511_), .Q(regs_23__9_) );
DFFPOSX1 DFFPOSX1_299 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_481_), .Q(regs_23__10_) );
DFFPOSX1 DFFPOSX1_300 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_482_), .Q(regs_23__11_) );
DFFPOSX1 DFFPOSX1_301 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_483_), .Q(regs_23__12_) );
DFFPOSX1 DFFPOSX1_302 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_484_), .Q(regs_23__13_) );
DFFPOSX1 DFFPOSX1_303 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_485_), .Q(regs_23__14_) );
DFFPOSX1 DFFPOSX1_304 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_486_), .Q(regs_23__15_) );
DFFPOSX1 DFFPOSX1_305 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_487_), .Q(regs_23__16_) );
DFFPOSX1 DFFPOSX1_306 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_488_), .Q(regs_23__17_) );
DFFPOSX1 DFFPOSX1_307 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_489_), .Q(regs_23__18_) );
DFFPOSX1 DFFPOSX1_308 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_490_), .Q(regs_23__19_) );
DFFPOSX1 DFFPOSX1_309 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_492_), .Q(regs_23__20_) );
DFFPOSX1 DFFPOSX1_310 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_493_), .Q(regs_23__21_) );
DFFPOSX1 DFFPOSX1_311 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_494_), .Q(regs_23__22_) );
DFFPOSX1 DFFPOSX1_312 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_495_), .Q(regs_23__23_) );
DFFPOSX1 DFFPOSX1_313 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_496_), .Q(regs_23__24_) );
DFFPOSX1 DFFPOSX1_314 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_497_), .Q(regs_23__25_) );
DFFPOSX1 DFFPOSX1_315 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_498_), .Q(regs_23__26_) );
DFFPOSX1 DFFPOSX1_316 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_499_), .Q(regs_23__27_) );
DFFPOSX1 DFFPOSX1_317 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_500_), .Q(regs_23__28_) );
DFFPOSX1 DFFPOSX1_318 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_501_), .Q(regs_23__29_) );
DFFPOSX1 DFFPOSX1_319 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_503_), .Q(regs_23__30_) );
DFFPOSX1 DFFPOSX1_320 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_504_), .Q(regs_23__31_) );
DFFPOSX1 DFFPOSX1_321 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_448_), .Q(regs_22__0_) );
DFFPOSX1 DFFPOSX1_322 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_459_), .Q(regs_22__1_) );
DFFPOSX1 DFFPOSX1_323 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_470_), .Q(regs_22__2_) );
DFFPOSX1 DFFPOSX1_324 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_473_), .Q(regs_22__3_) );
DFFPOSX1 DFFPOSX1_325 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_474_), .Q(regs_22__4_) );
DFFPOSX1 DFFPOSX1_326 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_475_), .Q(regs_22__5_) );
DFFPOSX1 DFFPOSX1_327 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_476_), .Q(regs_22__6_) );
DFFPOSX1 DFFPOSX1_328 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_477_), .Q(regs_22__7_) );
DFFPOSX1 DFFPOSX1_329 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_478_), .Q(regs_22__8_) );
DFFPOSX1 DFFPOSX1_330 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_479_), .Q(regs_22__9_) );
DFFPOSX1 DFFPOSX1_331 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_449_), .Q(regs_22__10_) );
DFFPOSX1 DFFPOSX1_332 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_450_), .Q(regs_22__11_) );
DFFPOSX1 DFFPOSX1_333 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_451_), .Q(regs_22__12_) );
DFFPOSX1 DFFPOSX1_334 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_452_), .Q(regs_22__13_) );
DFFPOSX1 DFFPOSX1_335 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_453_), .Q(regs_22__14_) );
DFFPOSX1 DFFPOSX1_336 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_454_), .Q(regs_22__15_) );
DFFPOSX1 DFFPOSX1_337 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_455_), .Q(regs_22__16_) );
DFFPOSX1 DFFPOSX1_338 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_456_), .Q(regs_22__17_) );
DFFPOSX1 DFFPOSX1_339 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_457_), .Q(regs_22__18_) );
DFFPOSX1 DFFPOSX1_340 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_458_), .Q(regs_22__19_) );
DFFPOSX1 DFFPOSX1_341 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_460_), .Q(regs_22__20_) );
DFFPOSX1 DFFPOSX1_342 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_461_), .Q(regs_22__21_) );
DFFPOSX1 DFFPOSX1_343 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_462_), .Q(regs_22__22_) );
DFFPOSX1 DFFPOSX1_344 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_463_), .Q(regs_22__23_) );
DFFPOSX1 DFFPOSX1_345 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_464_), .Q(regs_22__24_) );
DFFPOSX1 DFFPOSX1_346 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_465_), .Q(regs_22__25_) );
DFFPOSX1 DFFPOSX1_347 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_466_), .Q(regs_22__26_) );
DFFPOSX1 DFFPOSX1_348 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_467_), .Q(regs_22__27_) );
DFFPOSX1 DFFPOSX1_349 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_468_), .Q(regs_22__28_) );
DFFPOSX1 DFFPOSX1_350 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_469_), .Q(regs_22__29_) );
DFFPOSX1 DFFPOSX1_351 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_471_), .Q(regs_22__30_) );
DFFPOSX1 DFFPOSX1_352 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_472_), .Q(regs_22__31_) );
DFFPOSX1 DFFPOSX1_353 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_384_), .Q(regs_20__0_) );
DFFPOSX1 DFFPOSX1_354 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_395_), .Q(regs_20__1_) );
DFFPOSX1 DFFPOSX1_355 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_406_), .Q(regs_20__2_) );
DFFPOSX1 DFFPOSX1_356 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_409_), .Q(regs_20__3_) );
DFFPOSX1 DFFPOSX1_357 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_410_), .Q(regs_20__4_) );
DFFPOSX1 DFFPOSX1_358 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_411_), .Q(regs_20__5_) );
DFFPOSX1 DFFPOSX1_359 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_412_), .Q(regs_20__6_) );
DFFPOSX1 DFFPOSX1_360 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_413_), .Q(regs_20__7_) );
DFFPOSX1 DFFPOSX1_361 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_414_), .Q(regs_20__8_) );
DFFPOSX1 DFFPOSX1_362 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_415_), .Q(regs_20__9_) );
DFFPOSX1 DFFPOSX1_363 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_385_), .Q(regs_20__10_) );
DFFPOSX1 DFFPOSX1_364 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_386_), .Q(regs_20__11_) );
DFFPOSX1 DFFPOSX1_365 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_387_), .Q(regs_20__12_) );
DFFPOSX1 DFFPOSX1_366 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_388_), .Q(regs_20__13_) );
DFFPOSX1 DFFPOSX1_367 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_389_), .Q(regs_20__14_) );
DFFPOSX1 DFFPOSX1_368 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_390_), .Q(regs_20__15_) );
DFFPOSX1 DFFPOSX1_369 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_391_), .Q(regs_20__16_) );
DFFPOSX1 DFFPOSX1_370 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_392_), .Q(regs_20__17_) );
DFFPOSX1 DFFPOSX1_371 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_393_), .Q(regs_20__18_) );
DFFPOSX1 DFFPOSX1_372 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_394_), .Q(regs_20__19_) );
DFFPOSX1 DFFPOSX1_373 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_396_), .Q(regs_20__20_) );
DFFPOSX1 DFFPOSX1_374 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_397_), .Q(regs_20__21_) );
DFFPOSX1 DFFPOSX1_375 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_398_), .Q(regs_20__22_) );
DFFPOSX1 DFFPOSX1_376 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_399_), .Q(regs_20__23_) );
DFFPOSX1 DFFPOSX1_377 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_400_), .Q(regs_20__24_) );
DFFPOSX1 DFFPOSX1_378 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_401_), .Q(regs_20__25_) );
DFFPOSX1 DFFPOSX1_379 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_402_), .Q(regs_20__26_) );
DFFPOSX1 DFFPOSX1_380 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_403_), .Q(regs_20__27_) );
DFFPOSX1 DFFPOSX1_381 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_404_), .Q(regs_20__28_) );
DFFPOSX1 DFFPOSX1_382 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_405_), .Q(regs_20__29_) );
DFFPOSX1 DFFPOSX1_383 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_407_), .Q(regs_20__30_) );
DFFPOSX1 DFFPOSX1_384 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_408_), .Q(regs_20__31_) );
DFFPOSX1 DFFPOSX1_385 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_416_), .Q(regs_21__0_) );
DFFPOSX1 DFFPOSX1_386 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_427_), .Q(regs_21__1_) );
DFFPOSX1 DFFPOSX1_387 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_438_), .Q(regs_21__2_) );
DFFPOSX1 DFFPOSX1_388 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_441_), .Q(regs_21__3_) );
DFFPOSX1 DFFPOSX1_389 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_442_), .Q(regs_21__4_) );
DFFPOSX1 DFFPOSX1_390 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_443_), .Q(regs_21__5_) );
DFFPOSX1 DFFPOSX1_391 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_444_), .Q(regs_21__6_) );
DFFPOSX1 DFFPOSX1_392 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_445_), .Q(regs_21__7_) );
DFFPOSX1 DFFPOSX1_393 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_446_), .Q(regs_21__8_) );
DFFPOSX1 DFFPOSX1_394 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_447_), .Q(regs_21__9_) );
DFFPOSX1 DFFPOSX1_395 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_417_), .Q(regs_21__10_) );
DFFPOSX1 DFFPOSX1_396 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_418_), .Q(regs_21__11_) );
DFFPOSX1 DFFPOSX1_397 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_419_), .Q(regs_21__12_) );
DFFPOSX1 DFFPOSX1_398 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_420_), .Q(regs_21__13_) );
DFFPOSX1 DFFPOSX1_399 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_421_), .Q(regs_21__14_) );
DFFPOSX1 DFFPOSX1_400 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_422_), .Q(regs_21__15_) );
DFFPOSX1 DFFPOSX1_401 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_423_), .Q(regs_21__16_) );
DFFPOSX1 DFFPOSX1_402 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_424_), .Q(regs_21__17_) );
DFFPOSX1 DFFPOSX1_403 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_425_), .Q(regs_21__18_) );
DFFPOSX1 DFFPOSX1_404 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_426_), .Q(regs_21__19_) );
DFFPOSX1 DFFPOSX1_405 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_428_), .Q(regs_21__20_) );
DFFPOSX1 DFFPOSX1_406 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_429_), .Q(regs_21__21_) );
DFFPOSX1 DFFPOSX1_407 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_430_), .Q(regs_21__22_) );
DFFPOSX1 DFFPOSX1_408 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_431_), .Q(regs_21__23_) );
DFFPOSX1 DFFPOSX1_409 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_432_), .Q(regs_21__24_) );
DFFPOSX1 DFFPOSX1_410 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_433_), .Q(regs_21__25_) );
DFFPOSX1 DFFPOSX1_411 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_434_), .Q(regs_21__26_) );
DFFPOSX1 DFFPOSX1_412 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_435_), .Q(regs_21__27_) );
DFFPOSX1 DFFPOSX1_413 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_436_), .Q(regs_21__28_) );
DFFPOSX1 DFFPOSX1_414 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_437_), .Q(regs_21__29_) );
DFFPOSX1 DFFPOSX1_415 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_439_), .Q(regs_21__30_) );
DFFPOSX1 DFFPOSX1_416 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_440_), .Q(regs_21__31_) );
DFFPOSX1 DFFPOSX1_417 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_320_), .Q(regs_19__0_) );
DFFPOSX1 DFFPOSX1_418 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_331_), .Q(regs_19__1_) );
DFFPOSX1 DFFPOSX1_419 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_342_), .Q(regs_19__2_) );
DFFPOSX1 DFFPOSX1_420 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_345_), .Q(regs_19__3_) );
DFFPOSX1 DFFPOSX1_421 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_346_), .Q(regs_19__4_) );
DFFPOSX1 DFFPOSX1_422 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_347_), .Q(regs_19__5_) );
DFFPOSX1 DFFPOSX1_423 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_348_), .Q(regs_19__6_) );
DFFPOSX1 DFFPOSX1_424 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_349_), .Q(regs_19__7_) );
DFFPOSX1 DFFPOSX1_425 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_350_), .Q(regs_19__8_) );
DFFPOSX1 DFFPOSX1_426 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_351_), .Q(regs_19__9_) );
DFFPOSX1 DFFPOSX1_427 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_321_), .Q(regs_19__10_) );
DFFPOSX1 DFFPOSX1_428 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_322_), .Q(regs_19__11_) );
DFFPOSX1 DFFPOSX1_429 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_323_), .Q(regs_19__12_) );
DFFPOSX1 DFFPOSX1_430 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_324_), .Q(regs_19__13_) );
DFFPOSX1 DFFPOSX1_431 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_325_), .Q(regs_19__14_) );
DFFPOSX1 DFFPOSX1_432 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_326_), .Q(regs_19__15_) );
DFFPOSX1 DFFPOSX1_433 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_327_), .Q(regs_19__16_) );
DFFPOSX1 DFFPOSX1_434 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_328_), .Q(regs_19__17_) );
DFFPOSX1 DFFPOSX1_435 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_329_), .Q(regs_19__18_) );
DFFPOSX1 DFFPOSX1_436 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_330_), .Q(regs_19__19_) );
DFFPOSX1 DFFPOSX1_437 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_332_), .Q(regs_19__20_) );
DFFPOSX1 DFFPOSX1_438 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_333_), .Q(regs_19__21_) );
DFFPOSX1 DFFPOSX1_439 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_334_), .Q(regs_19__22_) );
DFFPOSX1 DFFPOSX1_440 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_335_), .Q(regs_19__23_) );
DFFPOSX1 DFFPOSX1_441 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_336_), .Q(regs_19__24_) );
DFFPOSX1 DFFPOSX1_442 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_337_), .Q(regs_19__25_) );
DFFPOSX1 DFFPOSX1_443 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_338_), .Q(regs_19__26_) );
DFFPOSX1 DFFPOSX1_444 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_339_), .Q(regs_19__27_) );
DFFPOSX1 DFFPOSX1_445 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_340_), .Q(regs_19__28_) );
DFFPOSX1 DFFPOSX1_446 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_341_), .Q(regs_19__29_) );
DFFPOSX1 DFFPOSX1_447 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_343_), .Q(regs_19__30_) );
DFFPOSX1 DFFPOSX1_448 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_344_), .Q(regs_19__31_) );
DFFPOSX1 DFFPOSX1_449 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_288_), .Q(regs_18__0_) );
DFFPOSX1 DFFPOSX1_450 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_299_), .Q(regs_18__1_) );
DFFPOSX1 DFFPOSX1_451 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_310_), .Q(regs_18__2_) );
DFFPOSX1 DFFPOSX1_452 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_313_), .Q(regs_18__3_) );
DFFPOSX1 DFFPOSX1_453 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_314_), .Q(regs_18__4_) );
DFFPOSX1 DFFPOSX1_454 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_315_), .Q(regs_18__5_) );
DFFPOSX1 DFFPOSX1_455 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_316_), .Q(regs_18__6_) );
DFFPOSX1 DFFPOSX1_456 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_317_), .Q(regs_18__7_) );
DFFPOSX1 DFFPOSX1_457 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_318_), .Q(regs_18__8_) );
DFFPOSX1 DFFPOSX1_458 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_319_), .Q(regs_18__9_) );
DFFPOSX1 DFFPOSX1_459 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_289_), .Q(regs_18__10_) );
DFFPOSX1 DFFPOSX1_460 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_290_), .Q(regs_18__11_) );
DFFPOSX1 DFFPOSX1_461 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_291_), .Q(regs_18__12_) );
DFFPOSX1 DFFPOSX1_462 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_292_), .Q(regs_18__13_) );
DFFPOSX1 DFFPOSX1_463 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_293_), .Q(regs_18__14_) );
DFFPOSX1 DFFPOSX1_464 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_294_), .Q(regs_18__15_) );
DFFPOSX1 DFFPOSX1_465 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_295_), .Q(regs_18__16_) );
DFFPOSX1 DFFPOSX1_466 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_296_), .Q(regs_18__17_) );
DFFPOSX1 DFFPOSX1_467 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_297_), .Q(regs_18__18_) );
DFFPOSX1 DFFPOSX1_468 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_298_), .Q(regs_18__19_) );
DFFPOSX1 DFFPOSX1_469 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_300_), .Q(regs_18__20_) );
DFFPOSX1 DFFPOSX1_470 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_301_), .Q(regs_18__21_) );
DFFPOSX1 DFFPOSX1_471 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_302_), .Q(regs_18__22_) );
DFFPOSX1 DFFPOSX1_472 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_303_), .Q(regs_18__23_) );
DFFPOSX1 DFFPOSX1_473 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_304_), .Q(regs_18__24_) );
DFFPOSX1 DFFPOSX1_474 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_305_), .Q(regs_18__25_) );
DFFPOSX1 DFFPOSX1_475 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_306_), .Q(regs_18__26_) );
DFFPOSX1 DFFPOSX1_476 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_307_), .Q(regs_18__27_) );
DFFPOSX1 DFFPOSX1_477 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_308_), .Q(regs_18__28_) );
DFFPOSX1 DFFPOSX1_478 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_309_), .Q(regs_18__29_) );
DFFPOSX1 DFFPOSX1_479 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_311_), .Q(regs_18__30_) );
DFFPOSX1 DFFPOSX1_480 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_312_), .Q(regs_18__31_) );
DFFPOSX1 DFFPOSX1_481 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_256_), .Q(regs_17__0_) );
DFFPOSX1 DFFPOSX1_482 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_267_), .Q(regs_17__1_) );
DFFPOSX1 DFFPOSX1_483 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_278_), .Q(regs_17__2_) );
DFFPOSX1 DFFPOSX1_484 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_281_), .Q(regs_17__3_) );
DFFPOSX1 DFFPOSX1_485 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_282_), .Q(regs_17__4_) );
DFFPOSX1 DFFPOSX1_486 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_283_), .Q(regs_17__5_) );
DFFPOSX1 DFFPOSX1_487 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_284_), .Q(regs_17__6_) );
DFFPOSX1 DFFPOSX1_488 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_285_), .Q(regs_17__7_) );
DFFPOSX1 DFFPOSX1_489 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_286_), .Q(regs_17__8_) );
DFFPOSX1 DFFPOSX1_490 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_287_), .Q(regs_17__9_) );
DFFPOSX1 DFFPOSX1_491 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_257_), .Q(regs_17__10_) );
DFFPOSX1 DFFPOSX1_492 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_258_), .Q(regs_17__11_) );
DFFPOSX1 DFFPOSX1_493 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_259_), .Q(regs_17__12_) );
DFFPOSX1 DFFPOSX1_494 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_260_), .Q(regs_17__13_) );
DFFPOSX1 DFFPOSX1_495 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_261_), .Q(regs_17__14_) );
DFFPOSX1 DFFPOSX1_496 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_262_), .Q(regs_17__15_) );
DFFPOSX1 DFFPOSX1_497 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_263_), .Q(regs_17__16_) );
DFFPOSX1 DFFPOSX1_498 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_264_), .Q(regs_17__17_) );
DFFPOSX1 DFFPOSX1_499 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_265_), .Q(regs_17__18_) );
DFFPOSX1 DFFPOSX1_500 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_266_), .Q(regs_17__19_) );
DFFPOSX1 DFFPOSX1_501 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_268_), .Q(regs_17__20_) );
DFFPOSX1 DFFPOSX1_502 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_269_), .Q(regs_17__21_) );
DFFPOSX1 DFFPOSX1_503 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_270_), .Q(regs_17__22_) );
DFFPOSX1 DFFPOSX1_504 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_271_), .Q(regs_17__23_) );
DFFPOSX1 DFFPOSX1_505 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_272_), .Q(regs_17__24_) );
DFFPOSX1 DFFPOSX1_506 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_273_), .Q(regs_17__25_) );
DFFPOSX1 DFFPOSX1_507 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_274_), .Q(regs_17__26_) );
DFFPOSX1 DFFPOSX1_508 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_275_), .Q(regs_17__27_) );
DFFPOSX1 DFFPOSX1_509 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_276_), .Q(regs_17__28_) );
DFFPOSX1 DFFPOSX1_510 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_277_), .Q(regs_17__29_) );
DFFPOSX1 DFFPOSX1_511 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_279_), .Q(regs_17__30_) );
DFFPOSX1 DFFPOSX1_512 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_280_), .Q(regs_17__31_) );
DFFPOSX1 DFFPOSX1_513 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_224_), .Q(regs_16__0_) );
DFFPOSX1 DFFPOSX1_514 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_235_), .Q(regs_16__1_) );
DFFPOSX1 DFFPOSX1_515 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_246_), .Q(regs_16__2_) );
DFFPOSX1 DFFPOSX1_516 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_249_), .Q(regs_16__3_) );
DFFPOSX1 DFFPOSX1_517 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_250_), .Q(regs_16__4_) );
DFFPOSX1 DFFPOSX1_518 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_251_), .Q(regs_16__5_) );
DFFPOSX1 DFFPOSX1_519 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_252_), .Q(regs_16__6_) );
DFFPOSX1 DFFPOSX1_520 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_253_), .Q(regs_16__7_) );
DFFPOSX1 DFFPOSX1_521 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_254_), .Q(regs_16__8_) );
DFFPOSX1 DFFPOSX1_522 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_255_), .Q(regs_16__9_) );
DFFPOSX1 DFFPOSX1_523 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_225_), .Q(regs_16__10_) );
DFFPOSX1 DFFPOSX1_524 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_226_), .Q(regs_16__11_) );
DFFPOSX1 DFFPOSX1_525 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_227_), .Q(regs_16__12_) );
DFFPOSX1 DFFPOSX1_526 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_228_), .Q(regs_16__13_) );
DFFPOSX1 DFFPOSX1_527 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_229_), .Q(regs_16__14_) );
DFFPOSX1 DFFPOSX1_528 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_230_), .Q(regs_16__15_) );
DFFPOSX1 DFFPOSX1_529 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_231_), .Q(regs_16__16_) );
DFFPOSX1 DFFPOSX1_530 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_232_), .Q(regs_16__17_) );
DFFPOSX1 DFFPOSX1_531 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_233_), .Q(regs_16__18_) );
DFFPOSX1 DFFPOSX1_532 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_234_), .Q(regs_16__19_) );
DFFPOSX1 DFFPOSX1_533 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_236_), .Q(regs_16__20_) );
DFFPOSX1 DFFPOSX1_534 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_237_), .Q(regs_16__21_) );
DFFPOSX1 DFFPOSX1_535 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_238_), .Q(regs_16__22_) );
DFFPOSX1 DFFPOSX1_536 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_239_), .Q(regs_16__23_) );
DFFPOSX1 DFFPOSX1_537 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_240_), .Q(regs_16__24_) );
DFFPOSX1 DFFPOSX1_538 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_241_), .Q(regs_16__25_) );
DFFPOSX1 DFFPOSX1_539 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_242_), .Q(regs_16__26_) );
DFFPOSX1 DFFPOSX1_540 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_243_), .Q(regs_16__27_) );
DFFPOSX1 DFFPOSX1_541 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_244_), .Q(regs_16__28_) );
DFFPOSX1 DFFPOSX1_542 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_245_), .Q(regs_16__29_) );
DFFPOSX1 DFFPOSX1_543 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_247_), .Q(regs_16__30_) );
DFFPOSX1 DFFPOSX1_544 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_248_), .Q(regs_16__31_) );
DFFPOSX1 DFFPOSX1_545 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_192_), .Q(regs_15__0_) );
DFFPOSX1 DFFPOSX1_546 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_203_), .Q(regs_15__1_) );
DFFPOSX1 DFFPOSX1_547 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_214_), .Q(regs_15__2_) );
DFFPOSX1 DFFPOSX1_548 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_217_), .Q(regs_15__3_) );
DFFPOSX1 DFFPOSX1_549 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_218_), .Q(regs_15__4_) );
DFFPOSX1 DFFPOSX1_550 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_219_), .Q(regs_15__5_) );
DFFPOSX1 DFFPOSX1_551 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_220_), .Q(regs_15__6_) );
DFFPOSX1 DFFPOSX1_552 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_221_), .Q(regs_15__7_) );
DFFPOSX1 DFFPOSX1_553 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_222_), .Q(regs_15__8_) );
DFFPOSX1 DFFPOSX1_554 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_223_), .Q(regs_15__9_) );
DFFPOSX1 DFFPOSX1_555 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_193_), .Q(regs_15__10_) );
DFFPOSX1 DFFPOSX1_556 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_194_), .Q(regs_15__11_) );
DFFPOSX1 DFFPOSX1_557 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_195_), .Q(regs_15__12_) );
DFFPOSX1 DFFPOSX1_558 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_196_), .Q(regs_15__13_) );
DFFPOSX1 DFFPOSX1_559 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_197_), .Q(regs_15__14_) );
DFFPOSX1 DFFPOSX1_560 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_198_), .Q(regs_15__15_) );
DFFPOSX1 DFFPOSX1_561 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_199_), .Q(regs_15__16_) );
DFFPOSX1 DFFPOSX1_562 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_200_), .Q(regs_15__17_) );
DFFPOSX1 DFFPOSX1_563 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_201_), .Q(regs_15__18_) );
DFFPOSX1 DFFPOSX1_564 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_202_), .Q(regs_15__19_) );
DFFPOSX1 DFFPOSX1_565 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_204_), .Q(regs_15__20_) );
DFFPOSX1 DFFPOSX1_566 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_205_), .Q(regs_15__21_) );
DFFPOSX1 DFFPOSX1_567 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_206_), .Q(regs_15__22_) );
DFFPOSX1 DFFPOSX1_568 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_207_), .Q(regs_15__23_) );
DFFPOSX1 DFFPOSX1_569 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_208_), .Q(regs_15__24_) );
DFFPOSX1 DFFPOSX1_570 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_209_), .Q(regs_15__25_) );
DFFPOSX1 DFFPOSX1_571 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_210_), .Q(regs_15__26_) );
DFFPOSX1 DFFPOSX1_572 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_211_), .Q(regs_15__27_) );
DFFPOSX1 DFFPOSX1_573 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_212_), .Q(regs_15__28_) );
DFFPOSX1 DFFPOSX1_574 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_213_), .Q(regs_15__29_) );
DFFPOSX1 DFFPOSX1_575 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_215_), .Q(regs_15__30_) );
DFFPOSX1 DFFPOSX1_576 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_216_), .Q(regs_15__31_) );
DFFPOSX1 DFFPOSX1_577 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_160_), .Q(regs_14__0_) );
DFFPOSX1 DFFPOSX1_578 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_171_), .Q(regs_14__1_) );
DFFPOSX1 DFFPOSX1_579 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_182_), .Q(regs_14__2_) );
DFFPOSX1 DFFPOSX1_580 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_185_), .Q(regs_14__3_) );
DFFPOSX1 DFFPOSX1_581 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_186_), .Q(regs_14__4_) );
DFFPOSX1 DFFPOSX1_582 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_187_), .Q(regs_14__5_) );
DFFPOSX1 DFFPOSX1_583 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_188_), .Q(regs_14__6_) );
DFFPOSX1 DFFPOSX1_584 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_189_), .Q(regs_14__7_) );
DFFPOSX1 DFFPOSX1_585 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_190_), .Q(regs_14__8_) );
DFFPOSX1 DFFPOSX1_586 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_191_), .Q(regs_14__9_) );
DFFPOSX1 DFFPOSX1_587 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_161_), .Q(regs_14__10_) );
DFFPOSX1 DFFPOSX1_588 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_162_), .Q(regs_14__11_) );
DFFPOSX1 DFFPOSX1_589 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_163_), .Q(regs_14__12_) );
DFFPOSX1 DFFPOSX1_590 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_164_), .Q(regs_14__13_) );
DFFPOSX1 DFFPOSX1_591 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_165_), .Q(regs_14__14_) );
DFFPOSX1 DFFPOSX1_592 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_166_), .Q(regs_14__15_) );
DFFPOSX1 DFFPOSX1_593 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_167_), .Q(regs_14__16_) );
DFFPOSX1 DFFPOSX1_594 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_168_), .Q(regs_14__17_) );
DFFPOSX1 DFFPOSX1_595 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_169_), .Q(regs_14__18_) );
DFFPOSX1 DFFPOSX1_596 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_170_), .Q(regs_14__19_) );
DFFPOSX1 DFFPOSX1_597 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_172_), .Q(regs_14__20_) );
DFFPOSX1 DFFPOSX1_598 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_173_), .Q(regs_14__21_) );
DFFPOSX1 DFFPOSX1_599 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_174_), .Q(regs_14__22_) );
DFFPOSX1 DFFPOSX1_600 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_175_), .Q(regs_14__23_) );
DFFPOSX1 DFFPOSX1_601 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_176_), .Q(regs_14__24_) );
DFFPOSX1 DFFPOSX1_602 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_177_), .Q(regs_14__25_) );
DFFPOSX1 DFFPOSX1_603 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_178_), .Q(regs_14__26_) );
DFFPOSX1 DFFPOSX1_604 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_179_), .Q(regs_14__27_) );
DFFPOSX1 DFFPOSX1_605 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_180_), .Q(regs_14__28_) );
DFFPOSX1 DFFPOSX1_606 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_181_), .Q(regs_14__29_) );
DFFPOSX1 DFFPOSX1_607 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_183_), .Q(regs_14__30_) );
DFFPOSX1 DFFPOSX1_608 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_184_), .Q(regs_14__31_) );
DFFPOSX1 DFFPOSX1_609 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_128_), .Q(regs_13__0_) );
DFFPOSX1 DFFPOSX1_610 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_139_), .Q(regs_13__1_) );
DFFPOSX1 DFFPOSX1_611 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_150_), .Q(regs_13__2_) );
DFFPOSX1 DFFPOSX1_612 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_153_), .Q(regs_13__3_) );
DFFPOSX1 DFFPOSX1_613 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_154_), .Q(regs_13__4_) );
DFFPOSX1 DFFPOSX1_614 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_155_), .Q(regs_13__5_) );
DFFPOSX1 DFFPOSX1_615 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_156_), .Q(regs_13__6_) );
DFFPOSX1 DFFPOSX1_616 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_157_), .Q(regs_13__7_) );
DFFPOSX1 DFFPOSX1_617 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_158_), .Q(regs_13__8_) );
DFFPOSX1 DFFPOSX1_618 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_159_), .Q(regs_13__9_) );
DFFPOSX1 DFFPOSX1_619 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_129_), .Q(regs_13__10_) );
DFFPOSX1 DFFPOSX1_620 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_130_), .Q(regs_13__11_) );
DFFPOSX1 DFFPOSX1_621 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_131_), .Q(regs_13__12_) );
DFFPOSX1 DFFPOSX1_622 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_132_), .Q(regs_13__13_) );
DFFPOSX1 DFFPOSX1_623 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_133_), .Q(regs_13__14_) );
DFFPOSX1 DFFPOSX1_624 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_134_), .Q(regs_13__15_) );
DFFPOSX1 DFFPOSX1_625 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_135_), .Q(regs_13__16_) );
DFFPOSX1 DFFPOSX1_626 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_136_), .Q(regs_13__17_) );
DFFPOSX1 DFFPOSX1_627 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_137_), .Q(regs_13__18_) );
DFFPOSX1 DFFPOSX1_628 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_138_), .Q(regs_13__19_) );
DFFPOSX1 DFFPOSX1_629 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_140_), .Q(regs_13__20_) );
DFFPOSX1 DFFPOSX1_630 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_141_), .Q(regs_13__21_) );
DFFPOSX1 DFFPOSX1_631 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_142_), .Q(regs_13__22_) );
DFFPOSX1 DFFPOSX1_632 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_143_), .Q(regs_13__23_) );
DFFPOSX1 DFFPOSX1_633 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_144_), .Q(regs_13__24_) );
DFFPOSX1 DFFPOSX1_634 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_145_), .Q(regs_13__25_) );
DFFPOSX1 DFFPOSX1_635 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_146_), .Q(regs_13__26_) );
DFFPOSX1 DFFPOSX1_636 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_147_), .Q(regs_13__27_) );
DFFPOSX1 DFFPOSX1_637 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_148_), .Q(regs_13__28_) );
DFFPOSX1 DFFPOSX1_638 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_149_), .Q(regs_13__29_) );
DFFPOSX1 DFFPOSX1_639 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_151_), .Q(regs_13__30_) );
DFFPOSX1 DFFPOSX1_640 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_152_), .Q(regs_13__31_) );
DFFPOSX1 DFFPOSX1_641 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_64_), .Q(regs_11__0_) );
DFFPOSX1 DFFPOSX1_642 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_75_), .Q(regs_11__1_) );
DFFPOSX1 DFFPOSX1_643 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_86_), .Q(regs_11__2_) );
DFFPOSX1 DFFPOSX1_644 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_89_), .Q(regs_11__3_) );
DFFPOSX1 DFFPOSX1_645 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_90_), .Q(regs_11__4_) );
DFFPOSX1 DFFPOSX1_646 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_91_), .Q(regs_11__5_) );
DFFPOSX1 DFFPOSX1_647 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_92_), .Q(regs_11__6_) );
DFFPOSX1 DFFPOSX1_648 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_93_), .Q(regs_11__7_) );
DFFPOSX1 DFFPOSX1_649 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_94_), .Q(regs_11__8_) );
DFFPOSX1 DFFPOSX1_650 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_95_), .Q(regs_11__9_) );
DFFPOSX1 DFFPOSX1_651 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_65_), .Q(regs_11__10_) );
DFFPOSX1 DFFPOSX1_652 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_66_), .Q(regs_11__11_) );
DFFPOSX1 DFFPOSX1_653 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_67_), .Q(regs_11__12_) );
DFFPOSX1 DFFPOSX1_654 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_68_), .Q(regs_11__13_) );
DFFPOSX1 DFFPOSX1_655 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_69_), .Q(regs_11__14_) );
DFFPOSX1 DFFPOSX1_656 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_70_), .Q(regs_11__15_) );
DFFPOSX1 DFFPOSX1_657 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_71_), .Q(regs_11__16_) );
DFFPOSX1 DFFPOSX1_658 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_72_), .Q(regs_11__17_) );
DFFPOSX1 DFFPOSX1_659 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_73_), .Q(regs_11__18_) );
DFFPOSX1 DFFPOSX1_660 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_74_), .Q(regs_11__19_) );
DFFPOSX1 DFFPOSX1_661 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_76_), .Q(regs_11__20_) );
DFFPOSX1 DFFPOSX1_662 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_77_), .Q(regs_11__21_) );
DFFPOSX1 DFFPOSX1_663 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_78_), .Q(regs_11__22_) );
DFFPOSX1 DFFPOSX1_664 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_79_), .Q(regs_11__23_) );
DFFPOSX1 DFFPOSX1_665 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_80_), .Q(regs_11__24_) );
DFFPOSX1 DFFPOSX1_666 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_81_), .Q(regs_11__25_) );
DFFPOSX1 DFFPOSX1_667 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_82_), .Q(regs_11__26_) );
DFFPOSX1 DFFPOSX1_668 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_83_), .Q(regs_11__27_) );
DFFPOSX1 DFFPOSX1_669 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_84_), .Q(regs_11__28_) );
DFFPOSX1 DFFPOSX1_670 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_85_), .Q(regs_11__29_) );
DFFPOSX1 DFFPOSX1_671 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_87_), .Q(regs_11__30_) );
DFFPOSX1 DFFPOSX1_672 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_88_), .Q(regs_11__31_) );
DFFPOSX1 DFFPOSX1_673 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_96_), .Q(regs_12__0_) );
DFFPOSX1 DFFPOSX1_674 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_107_), .Q(regs_12__1_) );
DFFPOSX1 DFFPOSX1_675 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_118_), .Q(regs_12__2_) );
DFFPOSX1 DFFPOSX1_676 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_121_), .Q(regs_12__3_) );
DFFPOSX1 DFFPOSX1_677 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_122_), .Q(regs_12__4_) );
DFFPOSX1 DFFPOSX1_678 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_123_), .Q(regs_12__5_) );
DFFPOSX1 DFFPOSX1_679 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_124_), .Q(regs_12__6_) );
DFFPOSX1 DFFPOSX1_680 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_125_), .Q(regs_12__7_) );
DFFPOSX1 DFFPOSX1_681 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_126_), .Q(regs_12__8_) );
DFFPOSX1 DFFPOSX1_682 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_127_), .Q(regs_12__9_) );
DFFPOSX1 DFFPOSX1_683 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_97_), .Q(regs_12__10_) );
DFFPOSX1 DFFPOSX1_684 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_98_), .Q(regs_12__11_) );
DFFPOSX1 DFFPOSX1_685 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_99_), .Q(regs_12__12_) );
DFFPOSX1 DFFPOSX1_686 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_100_), .Q(regs_12__13_) );
DFFPOSX1 DFFPOSX1_687 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_101_), .Q(regs_12__14_) );
DFFPOSX1 DFFPOSX1_688 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_102_), .Q(regs_12__15_) );
DFFPOSX1 DFFPOSX1_689 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_103_), .Q(regs_12__16_) );
DFFPOSX1 DFFPOSX1_690 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_104_), .Q(regs_12__17_) );
DFFPOSX1 DFFPOSX1_691 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_105_), .Q(regs_12__18_) );
DFFPOSX1 DFFPOSX1_692 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_106_), .Q(regs_12__19_) );
DFFPOSX1 DFFPOSX1_693 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_108_), .Q(regs_12__20_) );
DFFPOSX1 DFFPOSX1_694 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_109_), .Q(regs_12__21_) );
DFFPOSX1 DFFPOSX1_695 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_110_), .Q(regs_12__22_) );
DFFPOSX1 DFFPOSX1_696 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_111_), .Q(regs_12__23_) );
DFFPOSX1 DFFPOSX1_697 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_112_), .Q(regs_12__24_) );
DFFPOSX1 DFFPOSX1_698 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_113_), .Q(regs_12__25_) );
DFFPOSX1 DFFPOSX1_699 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_114_), .Q(regs_12__26_) );
DFFPOSX1 DFFPOSX1_700 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_115_), .Q(regs_12__27_) );
DFFPOSX1 DFFPOSX1_701 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_116_), .Q(regs_12__28_) );
DFFPOSX1 DFFPOSX1_702 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_117_), .Q(regs_12__29_) );
DFFPOSX1 DFFPOSX1_703 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_119_), .Q(regs_12__30_) );
DFFPOSX1 DFFPOSX1_704 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_120_), .Q(regs_12__31_) );
DFFPOSX1 DFFPOSX1_705 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_32_), .Q(regs_10__0_) );
DFFPOSX1 DFFPOSX1_706 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_43_), .Q(regs_10__1_) );
DFFPOSX1 DFFPOSX1_707 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_54_), .Q(regs_10__2_) );
DFFPOSX1 DFFPOSX1_708 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_57_), .Q(regs_10__3_) );
DFFPOSX1 DFFPOSX1_709 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_58_), .Q(regs_10__4_) );
DFFPOSX1 DFFPOSX1_710 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_59_), .Q(regs_10__5_) );
DFFPOSX1 DFFPOSX1_711 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_60_), .Q(regs_10__6_) );
DFFPOSX1 DFFPOSX1_712 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_61_), .Q(regs_10__7_) );
DFFPOSX1 DFFPOSX1_713 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_62_), .Q(regs_10__8_) );
DFFPOSX1 DFFPOSX1_714 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_63_), .Q(regs_10__9_) );
DFFPOSX1 DFFPOSX1_715 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_33_), .Q(regs_10__10_) );
DFFPOSX1 DFFPOSX1_716 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_34_), .Q(regs_10__11_) );
DFFPOSX1 DFFPOSX1_717 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_35_), .Q(regs_10__12_) );
DFFPOSX1 DFFPOSX1_718 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_36_), .Q(regs_10__13_) );
DFFPOSX1 DFFPOSX1_719 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_37_), .Q(regs_10__14_) );
DFFPOSX1 DFFPOSX1_720 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_38_), .Q(regs_10__15_) );
DFFPOSX1 DFFPOSX1_721 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_39_), .Q(regs_10__16_) );
DFFPOSX1 DFFPOSX1_722 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_40_), .Q(regs_10__17_) );
DFFPOSX1 DFFPOSX1_723 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_41_), .Q(regs_10__18_) );
DFFPOSX1 DFFPOSX1_724 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_42_), .Q(regs_10__19_) );
DFFPOSX1 DFFPOSX1_725 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_44_), .Q(regs_10__20_) );
DFFPOSX1 DFFPOSX1_726 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_45_), .Q(regs_10__21_) );
DFFPOSX1 DFFPOSX1_727 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_46_), .Q(regs_10__22_) );
DFFPOSX1 DFFPOSX1_728 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_47_), .Q(regs_10__23_) );
DFFPOSX1 DFFPOSX1_729 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_48_), .Q(regs_10__24_) );
DFFPOSX1 DFFPOSX1_730 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_49_), .Q(regs_10__25_) );
DFFPOSX1 DFFPOSX1_731 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_50_), .Q(regs_10__26_) );
DFFPOSX1 DFFPOSX1_732 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_51_), .Q(regs_10__27_) );
DFFPOSX1 DFFPOSX1_733 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_52_), .Q(regs_10__28_) );
DFFPOSX1 DFFPOSX1_734 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_53_), .Q(regs_10__29_) );
DFFPOSX1 DFFPOSX1_735 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_55_), .Q(regs_10__30_) );
DFFPOSX1 DFFPOSX1_736 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_56_), .Q(regs_10__31_) );
DFFPOSX1 DFFPOSX1_737 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_960_), .Q(regs_9__0_) );
DFFPOSX1 DFFPOSX1_738 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_971_), .Q(regs_9__1_) );
DFFPOSX1 DFFPOSX1_739 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_982_), .Q(regs_9__2_) );
DFFPOSX1 DFFPOSX1_740 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_985_), .Q(regs_9__3_) );
DFFPOSX1 DFFPOSX1_741 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_986_), .Q(regs_9__4_) );
DFFPOSX1 DFFPOSX1_742 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_987_), .Q(regs_9__5_) );
DFFPOSX1 DFFPOSX1_743 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_988_), .Q(regs_9__6_) );
DFFPOSX1 DFFPOSX1_744 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_989_), .Q(regs_9__7_) );
DFFPOSX1 DFFPOSX1_745 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_990_), .Q(regs_9__8_) );
DFFPOSX1 DFFPOSX1_746 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_991_), .Q(regs_9__9_) );
DFFPOSX1 DFFPOSX1_747 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_961_), .Q(regs_9__10_) );
DFFPOSX1 DFFPOSX1_748 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_962_), .Q(regs_9__11_) );
DFFPOSX1 DFFPOSX1_749 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_963_), .Q(regs_9__12_) );
DFFPOSX1 DFFPOSX1_750 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_964_), .Q(regs_9__13_) );
DFFPOSX1 DFFPOSX1_751 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_965_), .Q(regs_9__14_) );
DFFPOSX1 DFFPOSX1_752 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_966_), .Q(regs_9__15_) );
DFFPOSX1 DFFPOSX1_753 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_967_), .Q(regs_9__16_) );
DFFPOSX1 DFFPOSX1_754 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_968_), .Q(regs_9__17_) );
DFFPOSX1 DFFPOSX1_755 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_969_), .Q(regs_9__18_) );
DFFPOSX1 DFFPOSX1_756 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_970_), .Q(regs_9__19_) );
DFFPOSX1 DFFPOSX1_757 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_972_), .Q(regs_9__20_) );
DFFPOSX1 DFFPOSX1_758 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_973_), .Q(regs_9__21_) );
DFFPOSX1 DFFPOSX1_759 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_974_), .Q(regs_9__22_) );
DFFPOSX1 DFFPOSX1_760 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_975_), .Q(regs_9__23_) );
DFFPOSX1 DFFPOSX1_761 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_976_), .Q(regs_9__24_) );
DFFPOSX1 DFFPOSX1_762 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_977_), .Q(regs_9__25_) );
DFFPOSX1 DFFPOSX1_763 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_978_), .Q(regs_9__26_) );
DFFPOSX1 DFFPOSX1_764 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_979_), .Q(regs_9__27_) );
DFFPOSX1 DFFPOSX1_765 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_980_), .Q(regs_9__28_) );
DFFPOSX1 DFFPOSX1_766 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_981_), .Q(regs_9__29_) );
DFFPOSX1 DFFPOSX1_767 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_983_), .Q(regs_9__30_) );
DFFPOSX1 DFFPOSX1_768 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_984_), .Q(regs_9__31_) );
DFFPOSX1 DFFPOSX1_769 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_928_), .Q(regs_8__0_) );
DFFPOSX1 DFFPOSX1_770 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_939_), .Q(regs_8__1_) );
DFFPOSX1 DFFPOSX1_771 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_950_), .Q(regs_8__2_) );
DFFPOSX1 DFFPOSX1_772 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_953_), .Q(regs_8__3_) );
DFFPOSX1 DFFPOSX1_773 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_954_), .Q(regs_8__4_) );
DFFPOSX1 DFFPOSX1_774 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_955_), .Q(regs_8__5_) );
DFFPOSX1 DFFPOSX1_775 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_956_), .Q(regs_8__6_) );
DFFPOSX1 DFFPOSX1_776 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_957_), .Q(regs_8__7_) );
DFFPOSX1 DFFPOSX1_777 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_958_), .Q(regs_8__8_) );
DFFPOSX1 DFFPOSX1_778 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_959_), .Q(regs_8__9_) );
DFFPOSX1 DFFPOSX1_779 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_929_), .Q(regs_8__10_) );
DFFPOSX1 DFFPOSX1_780 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_930_), .Q(regs_8__11_) );
DFFPOSX1 DFFPOSX1_781 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_931_), .Q(regs_8__12_) );
DFFPOSX1 DFFPOSX1_782 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_932_), .Q(regs_8__13_) );
DFFPOSX1 DFFPOSX1_783 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_933_), .Q(regs_8__14_) );
DFFPOSX1 DFFPOSX1_784 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_934_), .Q(regs_8__15_) );
DFFPOSX1 DFFPOSX1_785 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_935_), .Q(regs_8__16_) );
DFFPOSX1 DFFPOSX1_786 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_936_), .Q(regs_8__17_) );
DFFPOSX1 DFFPOSX1_787 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_937_), .Q(regs_8__18_) );
DFFPOSX1 DFFPOSX1_788 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_938_), .Q(regs_8__19_) );
DFFPOSX1 DFFPOSX1_789 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_940_), .Q(regs_8__20_) );
DFFPOSX1 DFFPOSX1_790 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_941_), .Q(regs_8__21_) );
DFFPOSX1 DFFPOSX1_791 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_942_), .Q(regs_8__22_) );
DFFPOSX1 DFFPOSX1_792 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_943_), .Q(regs_8__23_) );
DFFPOSX1 DFFPOSX1_793 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_944_), .Q(regs_8__24_) );
DFFPOSX1 DFFPOSX1_794 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_945_), .Q(regs_8__25_) );
DFFPOSX1 DFFPOSX1_795 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_946_), .Q(regs_8__26_) );
DFFPOSX1 DFFPOSX1_796 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_947_), .Q(regs_8__27_) );
DFFPOSX1 DFFPOSX1_797 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_948_), .Q(regs_8__28_) );
DFFPOSX1 DFFPOSX1_798 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_949_), .Q(regs_8__29_) );
DFFPOSX1 DFFPOSX1_799 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_951_), .Q(regs_8__30_) );
DFFPOSX1 DFFPOSX1_800 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_952_), .Q(regs_8__31_) );
DFFPOSX1 DFFPOSX1_801 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_800_), .Q(regs_4__0_) );
DFFPOSX1 DFFPOSX1_802 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_811_), .Q(regs_4__1_) );
DFFPOSX1 DFFPOSX1_803 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_822_), .Q(regs_4__2_) );
DFFPOSX1 DFFPOSX1_804 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_825_), .Q(regs_4__3_) );
DFFPOSX1 DFFPOSX1_805 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_826_), .Q(regs_4__4_) );
DFFPOSX1 DFFPOSX1_806 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_827_), .Q(regs_4__5_) );
DFFPOSX1 DFFPOSX1_807 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_828_), .Q(regs_4__6_) );
DFFPOSX1 DFFPOSX1_808 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_829_), .Q(regs_4__7_) );
DFFPOSX1 DFFPOSX1_809 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_830_), .Q(regs_4__8_) );
DFFPOSX1 DFFPOSX1_810 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_831_), .Q(regs_4__9_) );
DFFPOSX1 DFFPOSX1_811 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_801_), .Q(regs_4__10_) );
DFFPOSX1 DFFPOSX1_812 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_802_), .Q(regs_4__11_) );
DFFPOSX1 DFFPOSX1_813 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_803_), .Q(regs_4__12_) );
DFFPOSX1 DFFPOSX1_814 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_804_), .Q(regs_4__13_) );
DFFPOSX1 DFFPOSX1_815 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_805_), .Q(regs_4__14_) );
DFFPOSX1 DFFPOSX1_816 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_806_), .Q(regs_4__15_) );
DFFPOSX1 DFFPOSX1_817 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_807_), .Q(regs_4__16_) );
DFFPOSX1 DFFPOSX1_818 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_808_), .Q(regs_4__17_) );
DFFPOSX1 DFFPOSX1_819 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_809_), .Q(regs_4__18_) );
DFFPOSX1 DFFPOSX1_820 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_810_), .Q(regs_4__19_) );
DFFPOSX1 DFFPOSX1_821 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_812_), .Q(regs_4__20_) );
DFFPOSX1 DFFPOSX1_822 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_813_), .Q(regs_4__21_) );
DFFPOSX1 DFFPOSX1_823 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_814_), .Q(regs_4__22_) );
DFFPOSX1 DFFPOSX1_824 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_815_), .Q(regs_4__23_) );
DFFPOSX1 DFFPOSX1_825 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_816_), .Q(regs_4__24_) );
DFFPOSX1 DFFPOSX1_826 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_817_), .Q(regs_4__25_) );
DFFPOSX1 DFFPOSX1_827 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_818_), .Q(regs_4__26_) );
DFFPOSX1 DFFPOSX1_828 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_819_), .Q(regs_4__27_) );
DFFPOSX1 DFFPOSX1_829 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_820_), .Q(regs_4__28_) );
DFFPOSX1 DFFPOSX1_830 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_821_), .Q(regs_4__29_) );
DFFPOSX1 DFFPOSX1_831 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_823_), .Q(regs_4__30_) );
DFFPOSX1 DFFPOSX1_832 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_824_), .Q(regs_4__31_) );
DFFPOSX1 DFFPOSX1_833 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_896_), .Q(regs_7__0_) );
DFFPOSX1 DFFPOSX1_834 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_907_), .Q(regs_7__1_) );
DFFPOSX1 DFFPOSX1_835 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_918_), .Q(regs_7__2_) );
DFFPOSX1 DFFPOSX1_836 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_921_), .Q(regs_7__3_) );
DFFPOSX1 DFFPOSX1_837 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_922_), .Q(regs_7__4_) );
DFFPOSX1 DFFPOSX1_838 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_923_), .Q(regs_7__5_) );
DFFPOSX1 DFFPOSX1_839 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_924_), .Q(regs_7__6_) );
DFFPOSX1 DFFPOSX1_840 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_925_), .Q(regs_7__7_) );
DFFPOSX1 DFFPOSX1_841 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_926_), .Q(regs_7__8_) );
DFFPOSX1 DFFPOSX1_842 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_927_), .Q(regs_7__9_) );
DFFPOSX1 DFFPOSX1_843 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_897_), .Q(regs_7__10_) );
DFFPOSX1 DFFPOSX1_844 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_898_), .Q(regs_7__11_) );
DFFPOSX1 DFFPOSX1_845 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_899_), .Q(regs_7__12_) );
DFFPOSX1 DFFPOSX1_846 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_900_), .Q(regs_7__13_) );
DFFPOSX1 DFFPOSX1_847 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_901_), .Q(regs_7__14_) );
DFFPOSX1 DFFPOSX1_848 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_902_), .Q(regs_7__15_) );
DFFPOSX1 DFFPOSX1_849 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_903_), .Q(regs_7__16_) );
DFFPOSX1 DFFPOSX1_850 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_904_), .Q(regs_7__17_) );
DFFPOSX1 DFFPOSX1_851 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_905_), .Q(regs_7__18_) );
DFFPOSX1 DFFPOSX1_852 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_906_), .Q(regs_7__19_) );
DFFPOSX1 DFFPOSX1_853 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_908_), .Q(regs_7__20_) );
DFFPOSX1 DFFPOSX1_854 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_909_), .Q(regs_7__21_) );
DFFPOSX1 DFFPOSX1_855 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_910_), .Q(regs_7__22_) );
DFFPOSX1 DFFPOSX1_856 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_911_), .Q(regs_7__23_) );
DFFPOSX1 DFFPOSX1_857 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_912_), .Q(regs_7__24_) );
DFFPOSX1 DFFPOSX1_858 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_913_), .Q(regs_7__25_) );
DFFPOSX1 DFFPOSX1_859 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_914_), .Q(regs_7__26_) );
DFFPOSX1 DFFPOSX1_860 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_915_), .Q(regs_7__27_) );
DFFPOSX1 DFFPOSX1_861 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_916_), .Q(regs_7__28_) );
DFFPOSX1 DFFPOSX1_862 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_917_), .Q(regs_7__29_) );
DFFPOSX1 DFFPOSX1_863 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_919_), .Q(regs_7__30_) );
DFFPOSX1 DFFPOSX1_864 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_920_), .Q(regs_7__31_) );
DFFPOSX1 DFFPOSX1_865 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_768_), .Q(regs_3__0_) );
DFFPOSX1 DFFPOSX1_866 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_779_), .Q(regs_3__1_) );
DFFPOSX1 DFFPOSX1_867 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_790_), .Q(regs_3__2_) );
DFFPOSX1 DFFPOSX1_868 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_793_), .Q(regs_3__3_) );
DFFPOSX1 DFFPOSX1_869 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_794_), .Q(regs_3__4_) );
DFFPOSX1 DFFPOSX1_870 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_795_), .Q(regs_3__5_) );
DFFPOSX1 DFFPOSX1_871 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_796_), .Q(regs_3__6_) );
DFFPOSX1 DFFPOSX1_872 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_797_), .Q(regs_3__7_) );
DFFPOSX1 DFFPOSX1_873 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_798_), .Q(regs_3__8_) );
DFFPOSX1 DFFPOSX1_874 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_799_), .Q(regs_3__9_) );
DFFPOSX1 DFFPOSX1_875 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_769_), .Q(regs_3__10_) );
DFFPOSX1 DFFPOSX1_876 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_770_), .Q(regs_3__11_) );
DFFPOSX1 DFFPOSX1_877 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_771_), .Q(regs_3__12_) );
DFFPOSX1 DFFPOSX1_878 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_772_), .Q(regs_3__13_) );
DFFPOSX1 DFFPOSX1_879 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_773_), .Q(regs_3__14_) );
DFFPOSX1 DFFPOSX1_880 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_774_), .Q(regs_3__15_) );
DFFPOSX1 DFFPOSX1_881 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_775_), .Q(regs_3__16_) );
DFFPOSX1 DFFPOSX1_882 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_776_), .Q(regs_3__17_) );
DFFPOSX1 DFFPOSX1_883 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_777_), .Q(regs_3__18_) );
DFFPOSX1 DFFPOSX1_884 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_778_), .Q(regs_3__19_) );
DFFPOSX1 DFFPOSX1_885 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_780_), .Q(regs_3__20_) );
DFFPOSX1 DFFPOSX1_886 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_781_), .Q(regs_3__21_) );
DFFPOSX1 DFFPOSX1_887 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_782_), .Q(regs_3__22_) );
DFFPOSX1 DFFPOSX1_888 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_783_), .Q(regs_3__23_) );
DFFPOSX1 DFFPOSX1_889 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_784_), .Q(regs_3__24_) );
DFFPOSX1 DFFPOSX1_890 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_785_), .Q(regs_3__25_) );
DFFPOSX1 DFFPOSX1_891 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_786_), .Q(regs_3__26_) );
DFFPOSX1 DFFPOSX1_892 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_787_), .Q(regs_3__27_) );
DFFPOSX1 DFFPOSX1_893 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_788_), .Q(regs_3__28_) );
DFFPOSX1 DFFPOSX1_894 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf96), .D(_789_), .Q(regs_3__29_) );
DFFPOSX1 DFFPOSX1_895 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf95), .D(_791_), .Q(regs_3__30_) );
DFFPOSX1 DFFPOSX1_896 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf94), .D(_792_), .Q(regs_3__31_) );
DFFPOSX1 DFFPOSX1_897 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf93), .D(_704_), .Q(regs_2__0_) );
DFFPOSX1 DFFPOSX1_898 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf92), .D(_715_), .Q(regs_2__1_) );
DFFPOSX1 DFFPOSX1_899 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf91), .D(_726_), .Q(regs_2__2_) );
DFFPOSX1 DFFPOSX1_900 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf90), .D(_729_), .Q(regs_2__3_) );
DFFPOSX1 DFFPOSX1_901 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf89), .D(_730_), .Q(regs_2__4_) );
DFFPOSX1 DFFPOSX1_902 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_731_), .Q(regs_2__5_) );
DFFPOSX1 DFFPOSX1_903 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_732_), .Q(regs_2__6_) );
DFFPOSX1 DFFPOSX1_904 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_733_), .Q(regs_2__7_) );
DFFPOSX1 DFFPOSX1_905 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_734_), .Q(regs_2__8_) );
DFFPOSX1 DFFPOSX1_906 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_735_), .Q(regs_2__9_) );
DFFPOSX1 DFFPOSX1_907 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_705_), .Q(regs_2__10_) );
DFFPOSX1 DFFPOSX1_908 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_706_), .Q(regs_2__11_) );
DFFPOSX1 DFFPOSX1_909 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_707_), .Q(regs_2__12_) );
DFFPOSX1 DFFPOSX1_910 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_708_), .Q(regs_2__13_) );
DFFPOSX1 DFFPOSX1_911 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_709_), .Q(regs_2__14_) );
DFFPOSX1 DFFPOSX1_912 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_710_), .Q(regs_2__15_) );
DFFPOSX1 DFFPOSX1_913 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_711_), .Q(regs_2__16_) );
DFFPOSX1 DFFPOSX1_914 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_712_), .Q(regs_2__17_) );
DFFPOSX1 DFFPOSX1_915 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_713_), .Q(regs_2__18_) );
DFFPOSX1 DFFPOSX1_916 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_714_), .Q(regs_2__19_) );
DFFPOSX1 DFFPOSX1_917 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_716_), .Q(regs_2__20_) );
DFFPOSX1 DFFPOSX1_918 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_717_), .Q(regs_2__21_) );
DFFPOSX1 DFFPOSX1_919 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_718_), .Q(regs_2__22_) );
DFFPOSX1 DFFPOSX1_920 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_719_), .Q(regs_2__23_) );
DFFPOSX1 DFFPOSX1_921 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_720_), .Q(regs_2__24_) );
DFFPOSX1 DFFPOSX1_922 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_721_), .Q(regs_2__25_) );
DFFPOSX1 DFFPOSX1_923 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_722_), .Q(regs_2__26_) );
DFFPOSX1 DFFPOSX1_924 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_723_), .Q(regs_2__27_) );
DFFPOSX1 DFFPOSX1_925 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_724_), .Q(regs_2__28_) );
DFFPOSX1 DFFPOSX1_926 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_725_), .Q(regs_2__29_) );
DFFPOSX1 DFFPOSX1_927 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_727_), .Q(regs_2__30_) );
DFFPOSX1 DFFPOSX1_928 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_728_), .Q(regs_2__31_) );
DFFPOSX1 DFFPOSX1_929 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_864_), .Q(regs_6__0_) );
DFFPOSX1 DFFPOSX1_930 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_875_), .Q(regs_6__1_) );
DFFPOSX1 DFFPOSX1_931 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_886_), .Q(regs_6__2_) );
DFFPOSX1 DFFPOSX1_932 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_889_), .Q(regs_6__3_) );
DFFPOSX1 DFFPOSX1_933 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_890_), .Q(regs_6__4_) );
DFFPOSX1 DFFPOSX1_934 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_891_), .Q(regs_6__5_) );
DFFPOSX1 DFFPOSX1_935 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_892_), .Q(regs_6__6_) );
DFFPOSX1 DFFPOSX1_936 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_893_), .Q(regs_6__7_) );
DFFPOSX1 DFFPOSX1_937 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_894_), .Q(regs_6__8_) );
DFFPOSX1 DFFPOSX1_938 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_895_), .Q(regs_6__9_) );
DFFPOSX1 DFFPOSX1_939 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_865_), .Q(regs_6__10_) );
DFFPOSX1 DFFPOSX1_940 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_866_), .Q(regs_6__11_) );
DFFPOSX1 DFFPOSX1_941 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_867_), .Q(regs_6__12_) );
DFFPOSX1 DFFPOSX1_942 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_868_), .Q(regs_6__13_) );
DFFPOSX1 DFFPOSX1_943 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_869_), .Q(regs_6__14_) );
DFFPOSX1 DFFPOSX1_944 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_870_), .Q(regs_6__15_) );
DFFPOSX1 DFFPOSX1_945 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_871_), .Q(regs_6__16_) );
DFFPOSX1 DFFPOSX1_946 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_872_), .Q(regs_6__17_) );
DFFPOSX1 DFFPOSX1_947 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_873_), .Q(regs_6__18_) );
DFFPOSX1 DFFPOSX1_948 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_874_), .Q(regs_6__19_) );
DFFPOSX1 DFFPOSX1_949 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_876_), .Q(regs_6__20_) );
DFFPOSX1 DFFPOSX1_950 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_877_), .Q(regs_6__21_) );
DFFPOSX1 DFFPOSX1_951 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_878_), .Q(regs_6__22_) );
DFFPOSX1 DFFPOSX1_952 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_879_), .Q(regs_6__23_) );
DFFPOSX1 DFFPOSX1_953 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_880_), .Q(regs_6__24_) );
DFFPOSX1 DFFPOSX1_954 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_881_), .Q(regs_6__25_) );
DFFPOSX1 DFFPOSX1_955 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_882_), .Q(regs_6__26_) );
DFFPOSX1 DFFPOSX1_956 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_883_), .Q(regs_6__27_) );
DFFPOSX1 DFFPOSX1_957 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_884_), .Q(regs_6__28_) );
DFFPOSX1 DFFPOSX1_958 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_885_), .Q(regs_6__29_) );
DFFPOSX1 DFFPOSX1_959 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_887_), .Q(regs_6__30_) );
DFFPOSX1 DFFPOSX1_960 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_888_), .Q(regs_6__31_) );
DFFPOSX1 DFFPOSX1_961 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_832_), .Q(regs_5__0_) );
DFFPOSX1 DFFPOSX1_962 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_843_), .Q(regs_5__1_) );
DFFPOSX1 DFFPOSX1_963 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_854_), .Q(regs_5__2_) );
DFFPOSX1 DFFPOSX1_964 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_857_), .Q(regs_5__3_) );
DFFPOSX1 DFFPOSX1_965 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_858_), .Q(regs_5__4_) );
DFFPOSX1 DFFPOSX1_966 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_859_), .Q(regs_5__5_) );
DFFPOSX1 DFFPOSX1_967 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_860_), .Q(regs_5__6_) );
DFFPOSX1 DFFPOSX1_968 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_861_), .Q(regs_5__7_) );
DFFPOSX1 DFFPOSX1_969 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_862_), .Q(regs_5__8_) );
DFFPOSX1 DFFPOSX1_970 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_863_), .Q(regs_5__9_) );
DFFPOSX1 DFFPOSX1_971 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_833_), .Q(regs_5__10_) );
DFFPOSX1 DFFPOSX1_972 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_834_), .Q(regs_5__11_) );
DFFPOSX1 DFFPOSX1_973 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_835_), .Q(regs_5__12_) );
DFFPOSX1 DFFPOSX1_974 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_836_), .Q(regs_5__13_) );
DFFPOSX1 DFFPOSX1_975 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_837_), .Q(regs_5__14_) );
DFFPOSX1 DFFPOSX1_976 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_838_), .Q(regs_5__15_) );
DFFPOSX1 DFFPOSX1_977 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_839_), .Q(regs_5__16_) );
DFFPOSX1 DFFPOSX1_978 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_840_), .Q(regs_5__17_) );
DFFPOSX1 DFFPOSX1_979 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_841_), .Q(regs_5__18_) );
DFFPOSX1 DFFPOSX1_980 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_842_), .Q(regs_5__19_) );
DFFPOSX1 DFFPOSX1_981 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_844_), .Q(regs_5__20_) );
DFFPOSX1 DFFPOSX1_982 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_845_), .Q(regs_5__21_) );
DFFPOSX1 DFFPOSX1_983 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_846_), .Q(regs_5__22_) );
DFFPOSX1 DFFPOSX1_984 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_847_), .Q(regs_5__23_) );
DFFPOSX1 DFFPOSX1_985 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_848_), .Q(regs_5__24_) );
DFFPOSX1 DFFPOSX1_986 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_849_), .Q(regs_5__25_) );
DFFPOSX1 DFFPOSX1_987 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_850_), .Q(regs_5__26_) );
DFFPOSX1 DFFPOSX1_988 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_851_), .Q(regs_5__27_) );
DFFPOSX1 DFFPOSX1_989 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_852_), .Q(regs_5__28_) );
DFFPOSX1 DFFPOSX1_990 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_853_), .Q(regs_5__29_) );
DFFPOSX1 DFFPOSX1_991 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf98), .D(_855_), .Q(regs_5__30_) );
DFFPOSX1 DFFPOSX1_992 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf97), .D(_856_), .Q(regs_5__31_) );
OAI21X1 OAI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_1936_), .B(_1902__bF_buf4), .C(_1937_), .Y(_72_) );
INVX2 INVX2_211 ( .gnd(gnd), .vdd(vdd), .A(regs_11__18_), .Y(_1938_) );
NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(wdata[18]), .B(_1902__bF_buf3), .Y(_1939_) );
OAI21X1 OAI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_1938_), .B(_1902__bF_buf2), .C(_1939_), .Y(_73_) );
INVX2 INVX2_212 ( .gnd(gnd), .vdd(vdd), .A(regs_11__19_), .Y(_1940_) );
NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(wdata[19]), .B(_1902__bF_buf1), .Y(_1941_) );
OAI21X1 OAI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_1940_), .B(_1902__bF_buf0), .C(_1941_), .Y(_74_) );
INVX2 INVX2_213 ( .gnd(gnd), .vdd(vdd), .A(regs_11__20_), .Y(_1942_) );
NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(wdata[20]), .B(_1902__bF_buf7), .Y(_1943_) );
OAI21X1 OAI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_1942_), .B(_1902__bF_buf6), .C(_1943_), .Y(_76_) );
INVX2 INVX2_214 ( .gnd(gnd), .vdd(vdd), .A(regs_11__21_), .Y(_1944_) );
NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(wdata[21]), .B(_1902__bF_buf5), .Y(_1945_) );
OAI21X1 OAI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_1944_), .B(_1902__bF_buf4), .C(_1945_), .Y(_77_) );
INVX2 INVX2_215 ( .gnd(gnd), .vdd(vdd), .A(regs_11__22_), .Y(_1946_) );
NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(wdata[22]), .B(_1902__bF_buf3), .Y(_1947_) );
OAI21X1 OAI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_1902__bF_buf2), .C(_1947_), .Y(_78_) );
INVX2 INVX2_216 ( .gnd(gnd), .vdd(vdd), .A(regs_11__23_), .Y(_1948_) );
NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(wdata[23]), .B(_1902__bF_buf1), .Y(_1949_) );
OAI21X1 OAI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_1948_), .B(_1902__bF_buf0), .C(_1949_), .Y(_79_) );
INVX2 INVX2_217 ( .gnd(gnd), .vdd(vdd), .A(regs_11__24_), .Y(_1950_) );
NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(wdata[24]), .B(_1902__bF_buf7), .Y(_1951_) );
OAI21X1 OAI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_1950_), .B(_1902__bF_buf6), .C(_1951_), .Y(_80_) );
INVX2 INVX2_218 ( .gnd(gnd), .vdd(vdd), .A(regs_11__25_), .Y(_1952_) );
NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(wdata[25]), .B(_1902__bF_buf5), .Y(_1953_) );
OAI21X1 OAI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_1952_), .B(_1902__bF_buf4), .C(_1953_), .Y(_81_) );
INVX2 INVX2_219 ( .gnd(gnd), .vdd(vdd), .A(regs_11__26_), .Y(_1954_) );
NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(wdata[26]), .B(_1902__bF_buf3), .Y(_1955_) );
OAI21X1 OAI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_1954_), .B(_1902__bF_buf2), .C(_1955_), .Y(_82_) );
INVX2 INVX2_220 ( .gnd(gnd), .vdd(vdd), .A(regs_11__27_), .Y(_1956_) );
NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(wdata[27]), .B(_1902__bF_buf1), .Y(_1957_) );
OAI21X1 OAI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_1956_), .B(_1902__bF_buf0), .C(_1957_), .Y(_83_) );
INVX2 INVX2_221 ( .gnd(gnd), .vdd(vdd), .A(regs_11__28_), .Y(_1958_) );
NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(wdata[28]), .B(_1902__bF_buf7), .Y(_1959_) );
OAI21X1 OAI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_1958_), .B(_1902__bF_buf6), .C(_1959_), .Y(_84_) );
INVX2 INVX2_222 ( .gnd(gnd), .vdd(vdd), .A(regs_11__29_), .Y(_1960_) );
NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(wdata[29]), .B(_1902__bF_buf5), .Y(_1961_) );
OAI21X1 OAI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_1960_), .B(_1902__bF_buf4), .C(_1961_), .Y(_85_) );
INVX2 INVX2_223 ( .gnd(gnd), .vdd(vdd), .A(regs_11__30_), .Y(_1962_) );
NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(wdata[30]), .B(_1902__bF_buf3), .Y(_1963_) );
OAI21X1 OAI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_1962_), .B(_1902__bF_buf2), .C(_1963_), .Y(_87_) );
INVX2 INVX2_224 ( .gnd(gnd), .vdd(vdd), .A(regs_11__31_), .Y(_1964_) );
NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(wdata[31]), .B(_1902__bF_buf1), .Y(_1965_) );
OAI21X1 OAI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_1964_), .B(_1902__bF_buf0), .C(_1965_), .Y(_88_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf6), .B(_1901__bF_buf4), .Y(_1966_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(regs_10__0_), .B(_1966__bF_buf7), .Y(_1967_) );
AOI21X1 AOI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_992__bF_buf1), .B(_1966__bF_buf6), .C(_1967_), .Y(_32_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(regs_10__1_), .B(_1966__bF_buf5), .Y(_1968_) );
AOI21X1 AOI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1003__bF_buf1), .B(_1966__bF_buf4), .C(_1968_), .Y(_43_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(regs_10__2_), .B(_1966__bF_buf3), .Y(_1969_) );
AOI21X1 AOI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf1), .B(_1966__bF_buf2), .C(_1969_), .Y(_54_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(regs_10__3_), .B(_1966__bF_buf1), .Y(_1970_) );
AOI21X1 AOI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1007__bF_buf1), .B(_1966__bF_buf0), .C(_1970_), .Y(_57_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(regs_10__4_), .B(_1966__bF_buf7), .Y(_1971_) );
AOI21X1 AOI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1009__bF_buf0), .B(_1966__bF_buf6), .C(_1971_), .Y(_58_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(regs_10__5_), .B(_1966__bF_buf5), .Y(_1972_) );
AOI21X1 AOI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1011__bF_buf0), .B(_1966__bF_buf4), .C(_1972_), .Y(_59_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(regs_10__6_), .B(_1966__bF_buf3), .Y(_1973_) );
AOI21X1 AOI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1013__bF_buf0), .B(_1966__bF_buf2), .C(_1973_), .Y(_60_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(regs_10__7_), .B(_1966__bF_buf1), .Y(_1974_) );
AOI21X1 AOI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1015__bF_buf0), .B(_1966__bF_buf0), .C(_1974_), .Y(_61_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(regs_10__8_), .B(_1966__bF_buf7), .Y(_1975_) );
AOI21X1 AOI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf0), .B(_1966__bF_buf6), .C(_1975_), .Y(_62_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(regs_10__9_), .B(_1966__bF_buf5), .Y(_1976_) );
AOI21X1 AOI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1019__bF_buf0), .B(_1966__bF_buf4), .C(_1976_), .Y(_63_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(regs_10__10_), .B(_1966__bF_buf3), .Y(_1977_) );
AOI21X1 AOI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1021__bF_buf0), .B(_1966__bF_buf2), .C(_1977_), .Y(_33_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(regs_10__11_), .B(_1966__bF_buf1), .Y(_1978_) );
AOI21X1 AOI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_1023__bF_buf0), .B(_1966__bF_buf0), .C(_1978_), .Y(_34_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(regs_10__12_), .B(_1966__bF_buf7), .Y(_1979_) );
AOI21X1 AOI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1025__bF_buf0), .B(_1966__bF_buf6), .C(_1979_), .Y(_35_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(regs_10__13_), .B(_1966__bF_buf5), .Y(_1980_) );
AOI21X1 AOI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1027__bF_buf0), .B(_1966__bF_buf4), .C(_1980_), .Y(_36_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(regs_10__14_), .B(_1966__bF_buf3), .Y(_1981_) );
AOI21X1 AOI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1029__bF_buf0), .B(_1966__bF_buf2), .C(_1981_), .Y(_37_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(regs_10__15_), .B(_1966__bF_buf1), .Y(_1982_) );
AOI21X1 AOI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf0), .B(_1966__bF_buf0), .C(_1982_), .Y(_38_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(regs_10__16_), .B(_1966__bF_buf7), .Y(_1983_) );
AOI21X1 AOI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1033__bF_buf0), .B(_1966__bF_buf6), .C(_1983_), .Y(_39_) );
NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(regs_10__17_), .B(_1966__bF_buf5), .Y(_1984_) );
AOI21X1 AOI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1035__bF_buf0), .B(_1966__bF_buf4), .C(_1984_), .Y(_40_) );
NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(regs_10__18_), .B(_1966__bF_buf3), .Y(_1985_) );
AOI21X1 AOI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_1037__bF_buf0), .B(_1966__bF_buf2), .C(_1985_), .Y(_41_) );
NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(regs_10__19_), .B(_1966__bF_buf1), .Y(_1986_) );
AOI21X1 AOI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1039__bF_buf0), .B(_1966__bF_buf0), .C(_1986_), .Y(_42_) );
NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(regs_10__20_), .B(_1966__bF_buf7), .Y(_1987_) );
AOI21X1 AOI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1041__bF_buf0), .B(_1966__bF_buf6), .C(_1987_), .Y(_44_) );
NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(regs_10__21_), .B(_1966__bF_buf5), .Y(_1988_) );
AOI21X1 AOI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1043__bF_buf0), .B(_1966__bF_buf4), .C(_1988_), .Y(_45_) );
NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(regs_10__22_), .B(_1966__bF_buf3), .Y(_1989_) );
AOI21X1 AOI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1045__bF_buf0), .B(_1966__bF_buf2), .C(_1989_), .Y(_46_) );
NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(regs_10__23_), .B(_1966__bF_buf1), .Y(_1990_) );
AOI21X1 AOI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1047__bF_buf0), .B(_1966__bF_buf0), .C(_1990_), .Y(_47_) );
NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(regs_10__24_), .B(_1966__bF_buf7), .Y(_1991_) );
AOI21X1 AOI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1049__bF_buf0), .B(_1966__bF_buf6), .C(_1991_), .Y(_48_) );
NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(regs_10__25_), .B(_1966__bF_buf5), .Y(_1992_) );
AOI21X1 AOI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1051__bF_buf0), .B(_1966__bF_buf4), .C(_1992_), .Y(_49_) );
NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(regs_10__26_), .B(_1966__bF_buf3), .Y(_1993_) );
AOI21X1 AOI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1053__bF_buf0), .B(_1966__bF_buf2), .C(_1993_), .Y(_50_) );
NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(regs_10__27_), .B(_1966__bF_buf1), .Y(_1994_) );
AOI21X1 AOI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1055__bF_buf0), .B(_1966__bF_buf0), .C(_1994_), .Y(_51_) );
NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(regs_10__28_), .B(_1966__bF_buf7), .Y(_1995_) );
AOI21X1 AOI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1057__bF_buf0), .B(_1966__bF_buf6), .C(_1995_), .Y(_52_) );
NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(regs_10__29_), .B(_1966__bF_buf5), .Y(_1996_) );
AOI21X1 AOI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1059__bF_buf0), .B(_1966__bF_buf4), .C(_1996_), .Y(_53_) );
NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(regs_10__30_), .B(_1966__bF_buf3), .Y(_1997_) );
AOI21X1 AOI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1061__bF_buf0), .B(_1966__bF_buf2), .C(_1997_), .Y(_55_) );
NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(regs_10__31_), .B(_1966__bF_buf1), .Y(_1998_) );
AOI21X1 AOI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1063__bF_buf0), .B(_1966__bF_buf0), .C(_1998_), .Y(_56_) );
INVX2 INVX2_225 ( .gnd(gnd), .vdd(vdd), .A(regs_9__0_), .Y(_1999_) );
NOR2X1 NOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf3), .B(_1070__bF_buf7), .Y(_2000_) );
NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(wdata[0]), .B(_2000__bF_buf7), .Y(_2001_) );
OAI21X1 OAI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_1999_), .B(_2000__bF_buf6), .C(_2001_), .Y(_960_) );
INVX2 INVX2_226 ( .gnd(gnd), .vdd(vdd), .A(regs_9__1_), .Y(_2002_) );
NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(wdata[1]), .B(_2000__bF_buf5), .Y(_2003_) );
OAI21X1 OAI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(_2002_), .B(_2000__bF_buf4), .C(_2003_), .Y(_971_) );
INVX2 INVX2_227 ( .gnd(gnd), .vdd(vdd), .A(regs_9__2_), .Y(_2004_) );
NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(wdata[2]), .B(_2000__bF_buf3), .Y(_2005_) );
OAI21X1 OAI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_2004_), .B(_2000__bF_buf2), .C(_2005_), .Y(_982_) );
INVX2 INVX2_228 ( .gnd(gnd), .vdd(vdd), .A(regs_9__3_), .Y(_2006_) );
NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(wdata[3]), .B(_2000__bF_buf1), .Y(_2007_) );
OAI21X1 OAI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .B(_2000__bF_buf0), .C(_2007_), .Y(_985_) );
INVX2 INVX2_229 ( .gnd(gnd), .vdd(vdd), .A(regs_9__4_), .Y(_2008_) );
NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(wdata[4]), .B(_2000__bF_buf7), .Y(_2009_) );
OAI21X1 OAI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(_2008_), .B(_2000__bF_buf6), .C(_2009_), .Y(_986_) );
INVX2 INVX2_230 ( .gnd(gnd), .vdd(vdd), .A(regs_9__5_), .Y(_2010_) );
NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(wdata[5]), .B(_2000__bF_buf5), .Y(_2011_) );
OAI21X1 OAI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(_2010_), .B(_2000__bF_buf4), .C(_2011_), .Y(_987_) );
INVX2 INVX2_231 ( .gnd(gnd), .vdd(vdd), .A(regs_9__6_), .Y(_2012_) );
NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(wdata[6]), .B(_2000__bF_buf3), .Y(_2013_) );
OAI21X1 OAI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(_2012_), .B(_2000__bF_buf2), .C(_2013_), .Y(_988_) );
INVX2 INVX2_232 ( .gnd(gnd), .vdd(vdd), .A(regs_9__7_), .Y(_2014_) );
NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(wdata[7]), .B(_2000__bF_buf1), .Y(_2015_) );
OAI21X1 OAI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(_2014_), .B(_2000__bF_buf0), .C(_2015_), .Y(_989_) );
INVX2 INVX2_233 ( .gnd(gnd), .vdd(vdd), .A(regs_9__8_), .Y(_2016_) );
NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(wdata[8]), .B(_2000__bF_buf7), .Y(_2017_) );
OAI21X1 OAI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_2016_), .B(_2000__bF_buf6), .C(_2017_), .Y(_990_) );
INVX2 INVX2_234 ( .gnd(gnd), .vdd(vdd), .A(regs_9__9_), .Y(_2018_) );
NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(wdata[9]), .B(_2000__bF_buf5), .Y(_2019_) );
OAI21X1 OAI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(_2018_), .B(_2000__bF_buf4), .C(_2019_), .Y(_991_) );
INVX2 INVX2_235 ( .gnd(gnd), .vdd(vdd), .A(regs_9__10_), .Y(_2020_) );
NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(wdata[10]), .B(_2000__bF_buf3), .Y(_2021_) );
OAI21X1 OAI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_2020_), .B(_2000__bF_buf2), .C(_2021_), .Y(_961_) );
INVX2 INVX2_236 ( .gnd(gnd), .vdd(vdd), .A(regs_9__11_), .Y(_2022_) );
NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(wdata[11]), .B(_2000__bF_buf1), .Y(_2023_) );
OAI21X1 OAI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(_2022_), .B(_2000__bF_buf0), .C(_2023_), .Y(_962_) );
INVX2 INVX2_237 ( .gnd(gnd), .vdd(vdd), .A(regs_9__12_), .Y(_2024_) );
NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(wdata[12]), .B(_2000__bF_buf7), .Y(_2025_) );
OAI21X1 OAI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(_2024_), .B(_2000__bF_buf6), .C(_2025_), .Y(_963_) );
INVX2 INVX2_238 ( .gnd(gnd), .vdd(vdd), .A(regs_9__13_), .Y(_2026_) );
NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(wdata[13]), .B(_2000__bF_buf5), .Y(_2027_) );
OAI21X1 OAI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_2026_), .B(_2000__bF_buf4), .C(_2027_), .Y(_964_) );
INVX2 INVX2_239 ( .gnd(gnd), .vdd(vdd), .A(regs_9__14_), .Y(_2028_) );
NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(wdata[14]), .B(_2000__bF_buf3), .Y(_2029_) );
OAI21X1 OAI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(_2028_), .B(_2000__bF_buf2), .C(_2029_), .Y(_965_) );
INVX2 INVX2_240 ( .gnd(gnd), .vdd(vdd), .A(regs_9__15_), .Y(_2030_) );
NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(wdata[15]), .B(_2000__bF_buf1), .Y(_2031_) );
OAI21X1 OAI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_2030_), .B(_2000__bF_buf0), .C(_2031_), .Y(_966_) );
INVX2 INVX2_241 ( .gnd(gnd), .vdd(vdd), .A(regs_9__16_), .Y(_2032_) );
NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(wdata[16]), .B(_2000__bF_buf7), .Y(_2033_) );
OAI21X1 OAI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(_2032_), .B(_2000__bF_buf6), .C(_2033_), .Y(_967_) );
INVX2 INVX2_242 ( .gnd(gnd), .vdd(vdd), .A(regs_9__17_), .Y(_2034_) );
NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(wdata[17]), .B(_2000__bF_buf5), .Y(_2035_) );
OAI21X1 OAI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(_2034_), .B(_2000__bF_buf4), .C(_2035_), .Y(_968_) );
INVX2 INVX2_243 ( .gnd(gnd), .vdd(vdd), .A(regs_9__18_), .Y(_2036_) );
NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(wdata[18]), .B(_2000__bF_buf3), .Y(_2037_) );
OAI21X1 OAI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_2036_), .B(_2000__bF_buf2), .C(_2037_), .Y(_969_) );
INVX2 INVX2_244 ( .gnd(gnd), .vdd(vdd), .A(regs_9__19_), .Y(_2038_) );
NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(wdata[19]), .B(_2000__bF_buf1), .Y(_2039_) );
OAI21X1 OAI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(_2038_), .B(_2000__bF_buf0), .C(_2039_), .Y(_970_) );
INVX2 INVX2_245 ( .gnd(gnd), .vdd(vdd), .A(regs_9__20_), .Y(_2040_) );
NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(wdata[20]), .B(_2000__bF_buf7), .Y(_2041_) );
OAI21X1 OAI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(_2040_), .B(_2000__bF_buf6), .C(_2041_), .Y(_972_) );
INVX2 INVX2_246 ( .gnd(gnd), .vdd(vdd), .A(regs_9__21_), .Y(_2042_) );
NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(wdata[21]), .B(_2000__bF_buf5), .Y(_2043_) );
OAI21X1 OAI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(_2042_), .B(_2000__bF_buf4), .C(_2043_), .Y(_973_) );
INVX2 INVX2_247 ( .gnd(gnd), .vdd(vdd), .A(regs_9__22_), .Y(_2044_) );
NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(wdata[22]), .B(_2000__bF_buf3), .Y(_2045_) );
OAI21X1 OAI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(_2044_), .B(_2000__bF_buf2), .C(_2045_), .Y(_974_) );
INVX2 INVX2_248 ( .gnd(gnd), .vdd(vdd), .A(regs_9__23_), .Y(_2046_) );
NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(wdata[23]), .B(_2000__bF_buf1), .Y(_2047_) );
OAI21X1 OAI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(_2046_), .B(_2000__bF_buf0), .C(_2047_), .Y(_975_) );
INVX2 INVX2_249 ( .gnd(gnd), .vdd(vdd), .A(regs_9__24_), .Y(_2048_) );
NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(wdata[24]), .B(_2000__bF_buf7), .Y(_2049_) );
OAI21X1 OAI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(_2048_), .B(_2000__bF_buf6), .C(_2049_), .Y(_976_) );
INVX2 INVX2_250 ( .gnd(gnd), .vdd(vdd), .A(regs_9__25_), .Y(_2050_) );
NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(wdata[25]), .B(_2000__bF_buf5), .Y(_2051_) );
OAI21X1 OAI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(_2050_), .B(_2000__bF_buf4), .C(_2051_), .Y(_977_) );
INVX2 INVX2_251 ( .gnd(gnd), .vdd(vdd), .A(regs_9__26_), .Y(_2052_) );
NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(wdata[26]), .B(_2000__bF_buf3), .Y(_2053_) );
OAI21X1 OAI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(_2052_), .B(_2000__bF_buf2), .C(_2053_), .Y(_978_) );
INVX2 INVX2_252 ( .gnd(gnd), .vdd(vdd), .A(regs_9__27_), .Y(_2054_) );
NAND2X1 NAND2X1_254 ( .gnd(gnd), .vdd(vdd), .A(wdata[27]), .B(_2000__bF_buf1), .Y(_2055_) );
OAI21X1 OAI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(_2054_), .B(_2000__bF_buf0), .C(_2055_), .Y(_979_) );
INVX2 INVX2_253 ( .gnd(gnd), .vdd(vdd), .A(regs_9__28_), .Y(_2056_) );
NAND2X1 NAND2X1_255 ( .gnd(gnd), .vdd(vdd), .A(wdata[28]), .B(_2000__bF_buf7), .Y(_2057_) );
OAI21X1 OAI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(_2056_), .B(_2000__bF_buf6), .C(_2057_), .Y(_980_) );
INVX2 INVX2_254 ( .gnd(gnd), .vdd(vdd), .A(regs_9__29_), .Y(_2058_) );
NAND2X1 NAND2X1_256 ( .gnd(gnd), .vdd(vdd), .A(wdata[29]), .B(_2000__bF_buf5), .Y(_2059_) );
OAI21X1 OAI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_2058_), .B(_2000__bF_buf4), .C(_2059_), .Y(_981_) );
INVX2 INVX2_255 ( .gnd(gnd), .vdd(vdd), .A(regs_9__30_), .Y(_2060_) );
NAND2X1 NAND2X1_257 ( .gnd(gnd), .vdd(vdd), .A(wdata[30]), .B(_2000__bF_buf3), .Y(_2061_) );
OAI21X1 OAI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(_2060_), .B(_2000__bF_buf2), .C(_2061_), .Y(_983_) );
INVX2 INVX2_256 ( .gnd(gnd), .vdd(vdd), .A(regs_9__31_), .Y(_2062_) );
NAND2X1 NAND2X1_258 ( .gnd(gnd), .vdd(vdd), .A(wdata[31]), .B(_2000__bF_buf1), .Y(_2063_) );
OAI21X1 OAI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(_2062_), .B(_2000__bF_buf0), .C(_2063_), .Y(_984_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf2), .B(_1104__bF_buf7), .Y(_2064_) );
OAI21X1 OAI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf1), .B(_1104__bF_buf6), .C(regs_8__0_), .Y(_2065_) );
OAI21X1 OAI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf4), .B(_992__bF_buf0), .C(_2065_), .Y(_928_) );
OAI21X1 OAI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf0), .B(_1104__bF_buf5), .C(regs_8__1_), .Y(_2066_) );
OAI21X1 OAI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf3), .B(_1003__bF_buf0), .C(_2066_), .Y(_939_) );
OAI21X1 OAI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf5), .B(_1104__bF_buf4), .C(regs_8__2_), .Y(_2067_) );
OAI21X1 OAI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf2), .B(_1005__bF_buf0), .C(_2067_), .Y(_950_) );
OAI21X1 OAI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf4), .B(_1104__bF_buf3), .C(regs_8__3_), .Y(_2068_) );
OAI21X1 OAI21X1_512 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf1), .B(_1007__bF_buf0), .C(_2068_), .Y(_953_) );
OAI21X1 OAI21X1_513 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf3), .B(_1104__bF_buf2), .C(regs_8__4_), .Y(_2069_) );
OAI21X1 OAI21X1_514 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf0), .B(_1009__bF_buf3), .C(_2069_), .Y(_954_) );
OAI21X1 OAI21X1_515 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf2), .B(_1104__bF_buf1), .C(regs_8__5_), .Y(_2070_) );
OAI21X1 OAI21X1_516 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf4), .B(_1011__bF_buf3), .C(_2070_), .Y(_955_) );
OAI21X1 OAI21X1_517 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf1), .B(_1104__bF_buf0), .C(regs_8__6_), .Y(_2071_) );
OAI21X1 OAI21X1_518 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf3), .B(_1013__bF_buf3), .C(_2071_), .Y(_956_) );
OAI21X1 OAI21X1_519 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf0), .B(_1104__bF_buf14), .C(regs_8__7_), .Y(_2072_) );
OAI21X1 OAI21X1_520 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf2), .B(_1015__bF_buf3), .C(_2072_), .Y(_957_) );
OAI21X1 OAI21X1_521 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf5), .B(_1104__bF_buf13), .C(regs_8__8_), .Y(_2073_) );
OAI21X1 OAI21X1_522 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf1), .B(_1017__bF_buf3), .C(_2073_), .Y(_958_) );
OAI21X1 OAI21X1_523 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf4), .B(_1104__bF_buf12), .C(regs_8__9_), .Y(_2074_) );
OAI21X1 OAI21X1_524 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf0), .B(_1019__bF_buf3), .C(_2074_), .Y(_959_) );
OAI21X1 OAI21X1_525 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf3), .B(_1104__bF_buf11), .C(regs_8__10_), .Y(_2075_) );
OAI21X1 OAI21X1_526 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf4), .B(_1021__bF_buf3), .C(_2075_), .Y(_929_) );
OAI21X1 OAI21X1_527 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf2), .B(_1104__bF_buf10), .C(regs_8__11_), .Y(_2076_) );
OAI21X1 OAI21X1_528 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf3), .B(_1023__bF_buf3), .C(_2076_), .Y(_930_) );
OAI21X1 OAI21X1_529 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf1), .B(_1104__bF_buf9), .C(regs_8__12_), .Y(_2077_) );
OAI21X1 OAI21X1_530 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf2), .B(_1025__bF_buf3), .C(_2077_), .Y(_931_) );
OAI21X1 OAI21X1_531 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf0), .B(_1104__bF_buf8), .C(regs_8__13_), .Y(_2078_) );
OAI21X1 OAI21X1_532 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf1), .B(_1027__bF_buf3), .C(_2078_), .Y(_932_) );
OAI21X1 OAI21X1_533 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf5), .B(_1104__bF_buf7), .C(regs_8__14_), .Y(_2079_) );
OAI21X1 OAI21X1_534 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf0), .B(_1029__bF_buf3), .C(_2079_), .Y(_933_) );
OAI21X1 OAI21X1_535 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf4), .B(_1104__bF_buf6), .C(regs_8__15_), .Y(_2080_) );
OAI21X1 OAI21X1_536 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf4), .B(_1031__bF_buf3), .C(_2080_), .Y(_934_) );
OAI21X1 OAI21X1_537 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf3), .B(_1104__bF_buf5), .C(regs_8__16_), .Y(_2081_) );
OAI21X1 OAI21X1_538 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf3), .B(_1033__bF_buf3), .C(_2081_), .Y(_935_) );
OAI21X1 OAI21X1_539 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf2), .B(_1104__bF_buf4), .C(regs_8__17_), .Y(_2082_) );
OAI21X1 OAI21X1_540 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf2), .B(_1035__bF_buf3), .C(_2082_), .Y(_936_) );
OAI21X1 OAI21X1_541 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf1), .B(_1104__bF_buf3), .C(regs_8__18_), .Y(_2083_) );
OAI21X1 OAI21X1_542 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf1), .B(_1037__bF_buf3), .C(_2083_), .Y(_937_) );
OAI21X1 OAI21X1_543 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf0), .B(_1104__bF_buf2), .C(regs_8__19_), .Y(_2084_) );
OAI21X1 OAI21X1_544 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf0), .B(_1039__bF_buf3), .C(_2084_), .Y(_938_) );
OAI21X1 OAI21X1_545 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf5), .B(_1104__bF_buf1), .C(regs_8__20_), .Y(_2085_) );
OAI21X1 OAI21X1_546 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf4), .B(_1041__bF_buf3), .C(_2085_), .Y(_940_) );
OAI21X1 OAI21X1_547 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf4), .B(_1104__bF_buf0), .C(regs_8__21_), .Y(_2086_) );
OAI21X1 OAI21X1_548 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf3), .B(_1043__bF_buf3), .C(_2086_), .Y(_941_) );
OAI21X1 OAI21X1_549 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf3), .B(_1104__bF_buf14), .C(regs_8__22_), .Y(_2087_) );
OAI21X1 OAI21X1_550 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf2), .B(_1045__bF_buf3), .C(_2087_), .Y(_942_) );
OAI21X1 OAI21X1_551 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf2), .B(_1104__bF_buf13), .C(regs_8__23_), .Y(_2088_) );
OAI21X1 OAI21X1_552 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf1), .B(_1047__bF_buf3), .C(_2088_), .Y(_943_) );
OAI21X1 OAI21X1_553 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf1), .B(_1104__bF_buf12), .C(regs_8__24_), .Y(_2089_) );
OAI21X1 OAI21X1_554 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf0), .B(_1049__bF_buf3), .C(_2089_), .Y(_944_) );
OAI21X1 OAI21X1_555 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf0), .B(_1104__bF_buf11), .C(regs_8__25_), .Y(_2090_) );
OAI21X1 OAI21X1_556 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf4), .B(_1051__bF_buf3), .C(_2090_), .Y(_945_) );
OAI21X1 OAI21X1_557 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf5), .B(_1104__bF_buf10), .C(regs_8__26_), .Y(_2091_) );
OAI21X1 OAI21X1_558 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf3), .B(_1053__bF_buf3), .C(_2091_), .Y(_946_) );
OAI21X1 OAI21X1_559 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf4), .B(_1104__bF_buf9), .C(regs_8__27_), .Y(_2092_) );
OAI21X1 OAI21X1_560 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf2), .B(_1055__bF_buf3), .C(_2092_), .Y(_947_) );
OAI21X1 OAI21X1_561 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf3), .B(_1104__bF_buf8), .C(regs_8__28_), .Y(_2093_) );
OAI21X1 OAI21X1_562 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf1), .B(_1057__bF_buf3), .C(_2093_), .Y(_948_) );
OAI21X1 OAI21X1_563 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf2), .B(_1104__bF_buf7), .C(regs_8__29_), .Y(_2094_) );
OAI21X1 OAI21X1_564 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf0), .B(_1059__bF_buf3), .C(_2094_), .Y(_949_) );
OAI21X1 OAI21X1_565 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf1), .B(_1104__bF_buf6), .C(regs_8__30_), .Y(_2095_) );
OAI21X1 OAI21X1_566 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf4), .B(_1061__bF_buf3), .C(_2095_), .Y(_951_) );
OAI21X1 OAI21X1_567 ( .gnd(gnd), .vdd(vdd), .A(_1901__bF_buf0), .B(_1104__bF_buf5), .C(regs_8__31_), .Y(_2096_) );
OAI21X1 OAI21X1_568 ( .gnd(gnd), .vdd(vdd), .A(_2064__bF_buf3), .B(_1063__bF_buf3), .C(_2096_), .Y(_952_) );
INVX2 INVX2_257 ( .gnd(gnd), .vdd(vdd), .A(regs_7__0_), .Y(_2097_) );
NAND2X1 NAND2X1_259 ( .gnd(gnd), .vdd(vdd), .A(waddr[4]), .B(waddr[3]), .Y(_2098_) );
NOR2X1 NOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(waddr[2]), .B(_2098_), .Y(_2099_) );
INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(_2099_), .Y(_2100_) );
NOR2X1 NOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1142__bF_buf1), .B(_2100__bF_buf8), .Y(_2101_) );
NAND2X1 NAND2X1_260 ( .gnd(gnd), .vdd(vdd), .A(wdata[0]), .B(_2101__bF_buf7), .Y(_2102_) );
OAI21X1 OAI21X1_569 ( .gnd(gnd), .vdd(vdd), .A(_2097_), .B(_2101__bF_buf6), .C(_2102_), .Y(_896_) );
INVX2 INVX2_258 ( .gnd(gnd), .vdd(vdd), .A(regs_7__1_), .Y(_2103_) );
NAND2X1 NAND2X1_261 ( .gnd(gnd), .vdd(vdd), .A(wdata[1]), .B(_2101__bF_buf5), .Y(_2104_) );
OAI21X1 OAI21X1_570 ( .gnd(gnd), .vdd(vdd), .A(_2103_), .B(_2101__bF_buf4), .C(_2104_), .Y(_907_) );
INVX2 INVX2_259 ( .gnd(gnd), .vdd(vdd), .A(regs_7__2_), .Y(_2105_) );
NAND2X1 NAND2X1_262 ( .gnd(gnd), .vdd(vdd), .A(wdata[2]), .B(_2101__bF_buf3), .Y(_2106_) );
OAI21X1 OAI21X1_571 ( .gnd(gnd), .vdd(vdd), .A(_2105_), .B(_2101__bF_buf2), .C(_2106_), .Y(_918_) );
INVX2 INVX2_260 ( .gnd(gnd), .vdd(vdd), .A(regs_7__3_), .Y(_2107_) );
NAND2X1 NAND2X1_263 ( .gnd(gnd), .vdd(vdd), .A(wdata[3]), .B(_2101__bF_buf1), .Y(_2108_) );
OAI21X1 OAI21X1_572 ( .gnd(gnd), .vdd(vdd), .A(_2107_), .B(_2101__bF_buf0), .C(_2108_), .Y(_921_) );
INVX2 INVX2_261 ( .gnd(gnd), .vdd(vdd), .A(regs_7__4_), .Y(_2109_) );
NAND2X1 NAND2X1_264 ( .gnd(gnd), .vdd(vdd), .A(wdata[4]), .B(_2101__bF_buf7), .Y(_2110_) );
OAI21X1 OAI21X1_573 ( .gnd(gnd), .vdd(vdd), .A(_2109_), .B(_2101__bF_buf6), .C(_2110_), .Y(_922_) );
INVX2 INVX2_262 ( .gnd(gnd), .vdd(vdd), .A(regs_7__5_), .Y(_2111_) );
NAND2X1 NAND2X1_265 ( .gnd(gnd), .vdd(vdd), .A(wdata[5]), .B(_2101__bF_buf5), .Y(_2112_) );
OAI21X1 OAI21X1_574 ( .gnd(gnd), .vdd(vdd), .A(_2111_), .B(_2101__bF_buf4), .C(_2112_), .Y(_923_) );
INVX2 INVX2_263 ( .gnd(gnd), .vdd(vdd), .A(regs_7__6_), .Y(_2113_) );
NAND2X1 NAND2X1_266 ( .gnd(gnd), .vdd(vdd), .A(wdata[6]), .B(_2101__bF_buf3), .Y(_2114_) );
OAI21X1 OAI21X1_575 ( .gnd(gnd), .vdd(vdd), .A(_2113_), .B(_2101__bF_buf2), .C(_2114_), .Y(_924_) );
INVX2 INVX2_264 ( .gnd(gnd), .vdd(vdd), .A(regs_7__7_), .Y(_2115_) );
NAND2X1 NAND2X1_267 ( .gnd(gnd), .vdd(vdd), .A(wdata[7]), .B(_2101__bF_buf1), .Y(_2116_) );
OAI21X1 OAI21X1_576 ( .gnd(gnd), .vdd(vdd), .A(_2115_), .B(_2101__bF_buf0), .C(_2116_), .Y(_925_) );
INVX2 INVX2_265 ( .gnd(gnd), .vdd(vdd), .A(regs_7__8_), .Y(_2117_) );
NAND2X1 NAND2X1_268 ( .gnd(gnd), .vdd(vdd), .A(wdata[8]), .B(_2101__bF_buf7), .Y(_2118_) );
OAI21X1 OAI21X1_577 ( .gnd(gnd), .vdd(vdd), .A(_2117_), .B(_2101__bF_buf6), .C(_2118_), .Y(_926_) );
INVX2 INVX2_266 ( .gnd(gnd), .vdd(vdd), .A(regs_7__9_), .Y(_2119_) );
NAND2X1 NAND2X1_269 ( .gnd(gnd), .vdd(vdd), .A(wdata[9]), .B(_2101__bF_buf5), .Y(_2120_) );
OAI21X1 OAI21X1_578 ( .gnd(gnd), .vdd(vdd), .A(_2119_), .B(_2101__bF_buf4), .C(_2120_), .Y(_927_) );
INVX2 INVX2_267 ( .gnd(gnd), .vdd(vdd), .A(regs_7__10_), .Y(_2121_) );
NAND2X1 NAND2X1_270 ( .gnd(gnd), .vdd(vdd), .A(wdata[10]), .B(_2101__bF_buf3), .Y(_2122_) );
OAI21X1 OAI21X1_579 ( .gnd(gnd), .vdd(vdd), .A(_2121_), .B(_2101__bF_buf2), .C(_2122_), .Y(_897_) );
INVX2 INVX2_268 ( .gnd(gnd), .vdd(vdd), .A(regs_7__11_), .Y(_2123_) );
NAND2X1 NAND2X1_271 ( .gnd(gnd), .vdd(vdd), .A(wdata[11]), .B(_2101__bF_buf1), .Y(_2124_) );
OAI21X1 OAI21X1_580 ( .gnd(gnd), .vdd(vdd), .A(_2123_), .B(_2101__bF_buf0), .C(_2124_), .Y(_898_) );
INVX2 INVX2_269 ( .gnd(gnd), .vdd(vdd), .A(regs_7__12_), .Y(_2125_) );
NAND2X1 NAND2X1_272 ( .gnd(gnd), .vdd(vdd), .A(wdata[12]), .B(_2101__bF_buf7), .Y(_2126_) );
OAI21X1 OAI21X1_581 ( .gnd(gnd), .vdd(vdd), .A(_2125_), .B(_2101__bF_buf6), .C(_2126_), .Y(_899_) );
INVX2 INVX2_270 ( .gnd(gnd), .vdd(vdd), .A(regs_7__13_), .Y(_2127_) );
NAND2X1 NAND2X1_273 ( .gnd(gnd), .vdd(vdd), .A(wdata[13]), .B(_2101__bF_buf5), .Y(_2128_) );
OAI21X1 OAI21X1_582 ( .gnd(gnd), .vdd(vdd), .A(_2127_), .B(_2101__bF_buf4), .C(_2128_), .Y(_900_) );
INVX2 INVX2_271 ( .gnd(gnd), .vdd(vdd), .A(regs_7__14_), .Y(_2129_) );
NAND2X1 NAND2X1_274 ( .gnd(gnd), .vdd(vdd), .A(wdata[14]), .B(_2101__bF_buf3), .Y(_2130_) );
OAI21X1 OAI21X1_583 ( .gnd(gnd), .vdd(vdd), .A(_2129_), .B(_2101__bF_buf2), .C(_2130_), .Y(_901_) );
INVX2 INVX2_272 ( .gnd(gnd), .vdd(vdd), .A(regs_7__15_), .Y(_2131_) );
NAND2X1 NAND2X1_275 ( .gnd(gnd), .vdd(vdd), .A(wdata[15]), .B(_2101__bF_buf1), .Y(_2132_) );
OAI21X1 OAI21X1_584 ( .gnd(gnd), .vdd(vdd), .A(_2131_), .B(_2101__bF_buf0), .C(_2132_), .Y(_902_) );
INVX2 INVX2_273 ( .gnd(gnd), .vdd(vdd), .A(regs_7__16_), .Y(_2133_) );
NAND2X1 NAND2X1_276 ( .gnd(gnd), .vdd(vdd), .A(wdata[16]), .B(_2101__bF_buf7), .Y(_2134_) );
OAI21X1 OAI21X1_585 ( .gnd(gnd), .vdd(vdd), .A(_2133_), .B(_2101__bF_buf6), .C(_2134_), .Y(_903_) );
INVX2 INVX2_274 ( .gnd(gnd), .vdd(vdd), .A(regs_7__17_), .Y(_2135_) );
NAND2X1 NAND2X1_277 ( .gnd(gnd), .vdd(vdd), .A(wdata[17]), .B(_2101__bF_buf5), .Y(_2136_) );
OAI21X1 OAI21X1_586 ( .gnd(gnd), .vdd(vdd), .A(_2135_), .B(_2101__bF_buf4), .C(_2136_), .Y(_904_) );
INVX2 INVX2_275 ( .gnd(gnd), .vdd(vdd), .A(regs_7__18_), .Y(_2137_) );
NAND2X1 NAND2X1_278 ( .gnd(gnd), .vdd(vdd), .A(wdata[18]), .B(_2101__bF_buf3), .Y(_2138_) );
OAI21X1 OAI21X1_587 ( .gnd(gnd), .vdd(vdd), .A(_2137_), .B(_2101__bF_buf2), .C(_2138_), .Y(_905_) );
INVX2 INVX2_276 ( .gnd(gnd), .vdd(vdd), .A(regs_7__19_), .Y(_2139_) );
NAND2X1 NAND2X1_279 ( .gnd(gnd), .vdd(vdd), .A(wdata[19]), .B(_2101__bF_buf1), .Y(_2140_) );
OAI21X1 OAI21X1_588 ( .gnd(gnd), .vdd(vdd), .A(_2139_), .B(_2101__bF_buf0), .C(_2140_), .Y(_906_) );
INVX2 INVX2_277 ( .gnd(gnd), .vdd(vdd), .A(regs_7__20_), .Y(_2141_) );
NAND2X1 NAND2X1_280 ( .gnd(gnd), .vdd(vdd), .A(wdata[20]), .B(_2101__bF_buf7), .Y(_2142_) );
OAI21X1 OAI21X1_589 ( .gnd(gnd), .vdd(vdd), .A(_2141_), .B(_2101__bF_buf6), .C(_2142_), .Y(_908_) );
INVX2 INVX2_278 ( .gnd(gnd), .vdd(vdd), .A(regs_7__21_), .Y(_2143_) );
NAND2X1 NAND2X1_281 ( .gnd(gnd), .vdd(vdd), .A(wdata[21]), .B(_2101__bF_buf5), .Y(_2144_) );
OAI21X1 OAI21X1_590 ( .gnd(gnd), .vdd(vdd), .A(_2143_), .B(_2101__bF_buf4), .C(_2144_), .Y(_909_) );
INVX2 INVX2_279 ( .gnd(gnd), .vdd(vdd), .A(regs_7__22_), .Y(_2145_) );
NAND2X1 NAND2X1_282 ( .gnd(gnd), .vdd(vdd), .A(wdata[22]), .B(_2101__bF_buf3), .Y(_2146_) );
OAI21X1 OAI21X1_591 ( .gnd(gnd), .vdd(vdd), .A(_2145_), .B(_2101__bF_buf2), .C(_2146_), .Y(_910_) );
INVX2 INVX2_280 ( .gnd(gnd), .vdd(vdd), .A(regs_7__23_), .Y(_2147_) );
NAND2X1 NAND2X1_283 ( .gnd(gnd), .vdd(vdd), .A(wdata[23]), .B(_2101__bF_buf1), .Y(_2148_) );
OAI21X1 OAI21X1_592 ( .gnd(gnd), .vdd(vdd), .A(_2147_), .B(_2101__bF_buf0), .C(_2148_), .Y(_911_) );
INVX2 INVX2_281 ( .gnd(gnd), .vdd(vdd), .A(regs_7__24_), .Y(_2149_) );
NAND2X1 NAND2X1_284 ( .gnd(gnd), .vdd(vdd), .A(wdata[24]), .B(_2101__bF_buf7), .Y(_2150_) );
OAI21X1 OAI21X1_593 ( .gnd(gnd), .vdd(vdd), .A(_2149_), .B(_2101__bF_buf6), .C(_2150_), .Y(_912_) );
INVX2 INVX2_282 ( .gnd(gnd), .vdd(vdd), .A(regs_7__25_), .Y(_2151_) );
NAND2X1 NAND2X1_285 ( .gnd(gnd), .vdd(vdd), .A(wdata[25]), .B(_2101__bF_buf5), .Y(_2152_) );
OAI21X1 OAI21X1_594 ( .gnd(gnd), .vdd(vdd), .A(_2151_), .B(_2101__bF_buf4), .C(_2152_), .Y(_913_) );
INVX2 INVX2_283 ( .gnd(gnd), .vdd(vdd), .A(regs_7__26_), .Y(_2153_) );
NAND2X1 NAND2X1_286 ( .gnd(gnd), .vdd(vdd), .A(wdata[26]), .B(_2101__bF_buf3), .Y(_2154_) );
OAI21X1 OAI21X1_595 ( .gnd(gnd), .vdd(vdd), .A(_2153_), .B(_2101__bF_buf2), .C(_2154_), .Y(_914_) );
INVX2 INVX2_284 ( .gnd(gnd), .vdd(vdd), .A(regs_7__27_), .Y(_2155_) );
NAND2X1 NAND2X1_287 ( .gnd(gnd), .vdd(vdd), .A(wdata[27]), .B(_2101__bF_buf1), .Y(_2156_) );
OAI21X1 OAI21X1_596 ( .gnd(gnd), .vdd(vdd), .A(_2155_), .B(_2101__bF_buf0), .C(_2156_), .Y(_915_) );
INVX2 INVX2_285 ( .gnd(gnd), .vdd(vdd), .A(regs_7__28_), .Y(_2157_) );
NAND2X1 NAND2X1_288 ( .gnd(gnd), .vdd(vdd), .A(wdata[28]), .B(_2101__bF_buf7), .Y(_2158_) );
OAI21X1 OAI21X1_597 ( .gnd(gnd), .vdd(vdd), .A(_2157_), .B(_2101__bF_buf6), .C(_2158_), .Y(_916_) );
INVX2 INVX2_286 ( .gnd(gnd), .vdd(vdd), .A(regs_7__29_), .Y(_2159_) );
NAND2X1 NAND2X1_289 ( .gnd(gnd), .vdd(vdd), .A(wdata[29]), .B(_2101__bF_buf5), .Y(_2160_) );
OAI21X1 OAI21X1_598 ( .gnd(gnd), .vdd(vdd), .A(_2159_), .B(_2101__bF_buf4), .C(_2160_), .Y(_917_) );
INVX2 INVX2_287 ( .gnd(gnd), .vdd(vdd), .A(regs_7__30_), .Y(_2161_) );
NAND2X1 NAND2X1_290 ( .gnd(gnd), .vdd(vdd), .A(wdata[30]), .B(_2101__bF_buf3), .Y(_2162_) );
OAI21X1 OAI21X1_599 ( .gnd(gnd), .vdd(vdd), .A(_2161_), .B(_2101__bF_buf2), .C(_2162_), .Y(_919_) );
INVX2 INVX2_288 ( .gnd(gnd), .vdd(vdd), .A(regs_7__31_), .Y(_2163_) );
NAND2X1 NAND2X1_291 ( .gnd(gnd), .vdd(vdd), .A(wdata[31]), .B(_2101__bF_buf1), .Y(_2164_) );
OAI21X1 OAI21X1_600 ( .gnd(gnd), .vdd(vdd), .A(_2163_), .B(_2101__bF_buf0), .C(_2164_), .Y(_920_) );
NAND2X1 NAND2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_998_), .B(_2099_), .Y(_2165_) );
OAI21X1 OAI21X1_601 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf5), .B(_2100__bF_buf7), .C(regs_6__0_), .Y(_2166_) );
OAI21X1 OAI21X1_602 ( .gnd(gnd), .vdd(vdd), .A(_992__bF_buf3), .B(_2165__bF_buf4), .C(_2166_), .Y(_864_) );
OAI21X1 OAI21X1_603 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf4), .B(_2100__bF_buf6), .C(regs_6__1_), .Y(_2167_) );
OAI21X1 OAI21X1_604 ( .gnd(gnd), .vdd(vdd), .A(_1003__bF_buf3), .B(_2165__bF_buf3), .C(_2167_), .Y(_875_) );
OAI21X1 OAI21X1_605 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf3), .B(_2100__bF_buf5), .C(regs_6__2_), .Y(_2168_) );
OAI21X1 OAI21X1_606 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf3), .B(_2165__bF_buf2), .C(_2168_), .Y(_886_) );
OAI21X1 OAI21X1_607 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf2), .B(_2100__bF_buf4), .C(regs_6__3_), .Y(_2169_) );
OAI21X1 OAI21X1_608 ( .gnd(gnd), .vdd(vdd), .A(_1007__bF_buf3), .B(_2165__bF_buf1), .C(_2169_), .Y(_889_) );
OAI21X1 OAI21X1_609 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf1), .B(_2100__bF_buf3), .C(regs_6__4_), .Y(_2170_) );
OAI21X1 OAI21X1_610 ( .gnd(gnd), .vdd(vdd), .A(_1009__bF_buf2), .B(_2165__bF_buf0), .C(_2170_), .Y(_890_) );
OAI21X1 OAI21X1_611 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf0), .B(_2100__bF_buf2), .C(regs_6__5_), .Y(_2171_) );
OAI21X1 OAI21X1_612 ( .gnd(gnd), .vdd(vdd), .A(_1011__bF_buf2), .B(_2165__bF_buf4), .C(_2171_), .Y(_891_) );
OAI21X1 OAI21X1_613 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf9), .B(_2100__bF_buf1), .C(regs_6__6_), .Y(_2172_) );
OAI21X1 OAI21X1_614 ( .gnd(gnd), .vdd(vdd), .A(_1013__bF_buf2), .B(_2165__bF_buf3), .C(_2172_), .Y(_892_) );
OAI21X1 OAI21X1_615 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf8), .B(_2100__bF_buf0), .C(regs_6__7_), .Y(_2173_) );
OAI21X1 OAI21X1_616 ( .gnd(gnd), .vdd(vdd), .A(_1015__bF_buf2), .B(_2165__bF_buf2), .C(_2173_), .Y(_893_) );
OAI21X1 OAI21X1_617 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf7), .B(_2100__bF_buf8), .C(regs_6__8_), .Y(_2174_) );
OAI21X1 OAI21X1_618 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf2), .B(_2165__bF_buf1), .C(_2174_), .Y(_894_) );
OAI21X1 OAI21X1_619 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf6), .B(_2100__bF_buf7), .C(regs_6__9_), .Y(_2175_) );
OAI21X1 OAI21X1_620 ( .gnd(gnd), .vdd(vdd), .A(_1019__bF_buf2), .B(_2165__bF_buf0), .C(_2175_), .Y(_895_) );
OAI21X1 OAI21X1_621 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf5), .B(_2100__bF_buf6), .C(regs_6__10_), .Y(_2176_) );
OAI21X1 OAI21X1_622 ( .gnd(gnd), .vdd(vdd), .A(_1021__bF_buf2), .B(_2165__bF_buf4), .C(_2176_), .Y(_865_) );
OAI21X1 OAI21X1_623 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf4), .B(_2100__bF_buf5), .C(regs_6__11_), .Y(_2177_) );
OAI21X1 OAI21X1_624 ( .gnd(gnd), .vdd(vdd), .A(_1023__bF_buf2), .B(_2165__bF_buf3), .C(_2177_), .Y(_866_) );
OAI21X1 OAI21X1_625 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf3), .B(_2100__bF_buf4), .C(regs_6__12_), .Y(_2178_) );
OAI21X1 OAI21X1_626 ( .gnd(gnd), .vdd(vdd), .A(_1025__bF_buf2), .B(_2165__bF_buf2), .C(_2178_), .Y(_867_) );
OAI21X1 OAI21X1_627 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf2), .B(_2100__bF_buf3), .C(regs_6__13_), .Y(_2179_) );
OAI21X1 OAI21X1_628 ( .gnd(gnd), .vdd(vdd), .A(_1027__bF_buf2), .B(_2165__bF_buf1), .C(_2179_), .Y(_868_) );
OAI21X1 OAI21X1_629 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf1), .B(_2100__bF_buf2), .C(regs_6__14_), .Y(_2180_) );
OAI21X1 OAI21X1_630 ( .gnd(gnd), .vdd(vdd), .A(_1029__bF_buf2), .B(_2165__bF_buf0), .C(_2180_), .Y(_869_) );
OAI21X1 OAI21X1_631 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf0), .B(_2100__bF_buf1), .C(regs_6__15_), .Y(_2181_) );
OAI21X1 OAI21X1_632 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf2), .B(_2165__bF_buf4), .C(_2181_), .Y(_870_) );
OAI21X1 OAI21X1_633 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf9), .B(_2100__bF_buf0), .C(regs_6__16_), .Y(_2182_) );
OAI21X1 OAI21X1_634 ( .gnd(gnd), .vdd(vdd), .A(_1033__bF_buf2), .B(_2165__bF_buf3), .C(_2182_), .Y(_871_) );
OAI21X1 OAI21X1_635 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf8), .B(_2100__bF_buf8), .C(regs_6__17_), .Y(_2183_) );
OAI21X1 OAI21X1_636 ( .gnd(gnd), .vdd(vdd), .A(_1035__bF_buf2), .B(_2165__bF_buf2), .C(_2183_), .Y(_872_) );
OAI21X1 OAI21X1_637 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf7), .B(_2100__bF_buf7), .C(regs_6__18_), .Y(_2184_) );
OAI21X1 OAI21X1_638 ( .gnd(gnd), .vdd(vdd), .A(_1037__bF_buf2), .B(_2165__bF_buf1), .C(_2184_), .Y(_873_) );
OAI21X1 OAI21X1_639 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf6), .B(_2100__bF_buf6), .C(regs_6__19_), .Y(_2185_) );
OAI21X1 OAI21X1_640 ( .gnd(gnd), .vdd(vdd), .A(_1039__bF_buf2), .B(_2165__bF_buf0), .C(_2185_), .Y(_874_) );
OAI21X1 OAI21X1_641 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf5), .B(_2100__bF_buf5), .C(regs_6__20_), .Y(_2186_) );
OAI21X1 OAI21X1_642 ( .gnd(gnd), .vdd(vdd), .A(_1041__bF_buf2), .B(_2165__bF_buf4), .C(_2186_), .Y(_876_) );
OAI21X1 OAI21X1_643 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf4), .B(_2100__bF_buf4), .C(regs_6__21_), .Y(_2187_) );
OAI21X1 OAI21X1_644 ( .gnd(gnd), .vdd(vdd), .A(_1043__bF_buf2), .B(_2165__bF_buf3), .C(_2187_), .Y(_877_) );
OAI21X1 OAI21X1_645 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf3), .B(_2100__bF_buf3), .C(regs_6__22_), .Y(_2188_) );
OAI21X1 OAI21X1_646 ( .gnd(gnd), .vdd(vdd), .A(_1045__bF_buf2), .B(_2165__bF_buf2), .C(_2188_), .Y(_878_) );
OAI21X1 OAI21X1_647 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf2), .B(_2100__bF_buf2), .C(regs_6__23_), .Y(_2189_) );
OAI21X1 OAI21X1_648 ( .gnd(gnd), .vdd(vdd), .A(_1047__bF_buf2), .B(_2165__bF_buf1), .C(_2189_), .Y(_879_) );
OAI21X1 OAI21X1_649 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf1), .B(_2100__bF_buf1), .C(regs_6__24_), .Y(_2190_) );
OAI21X1 OAI21X1_650 ( .gnd(gnd), .vdd(vdd), .A(_1049__bF_buf2), .B(_2165__bF_buf0), .C(_2190_), .Y(_880_) );
OAI21X1 OAI21X1_651 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf0), .B(_2100__bF_buf0), .C(regs_6__25_), .Y(_2191_) );
OAI21X1 OAI21X1_652 ( .gnd(gnd), .vdd(vdd), .A(_1051__bF_buf2), .B(_2165__bF_buf4), .C(_2191_), .Y(_881_) );
OAI21X1 OAI21X1_653 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf9), .B(_2100__bF_buf8), .C(regs_6__26_), .Y(_2192_) );
OAI21X1 OAI21X1_654 ( .gnd(gnd), .vdd(vdd), .A(_1053__bF_buf2), .B(_2165__bF_buf3), .C(_2192_), .Y(_882_) );
OAI21X1 OAI21X1_655 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf8), .B(_2100__bF_buf7), .C(regs_6__27_), .Y(_2193_) );
OAI21X1 OAI21X1_656 ( .gnd(gnd), .vdd(vdd), .A(_1055__bF_buf2), .B(_2165__bF_buf2), .C(_2193_), .Y(_883_) );
OAI21X1 OAI21X1_657 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf7), .B(_2100__bF_buf6), .C(regs_6__28_), .Y(_2194_) );
OAI21X1 OAI21X1_658 ( .gnd(gnd), .vdd(vdd), .A(_1057__bF_buf2), .B(_2165__bF_buf1), .C(_2194_), .Y(_884_) );
OAI21X1 OAI21X1_659 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf6), .B(_2100__bF_buf5), .C(regs_6__29_), .Y(_2195_) );
OAI21X1 OAI21X1_660 ( .gnd(gnd), .vdd(vdd), .A(_1059__bF_buf2), .B(_2165__bF_buf0), .C(_2195_), .Y(_885_) );
OAI21X1 OAI21X1_661 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf5), .B(_2100__bF_buf4), .C(regs_6__30_), .Y(_2196_) );
OAI21X1 OAI21X1_662 ( .gnd(gnd), .vdd(vdd), .A(_1061__bF_buf2), .B(_2165__bF_buf4), .C(_2196_), .Y(_887_) );
OAI21X1 OAI21X1_663 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf4), .B(_2100__bF_buf3), .C(regs_6__31_), .Y(_2197_) );
OAI21X1 OAI21X1_664 ( .gnd(gnd), .vdd(vdd), .A(_1063__bF_buf2), .B(_2165__bF_buf3), .C(_2197_), .Y(_888_) );
NAND2X1 NAND2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_2099_), .B(_1068_), .Y(_2198_) );
OAI21X1 OAI21X1_665 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf6), .B(_2100__bF_buf2), .C(regs_5__0_), .Y(_2199_) );
OAI21X1 OAI21X1_666 ( .gnd(gnd), .vdd(vdd), .A(_992__bF_buf2), .B(_2198__bF_buf4), .C(_2199_), .Y(_832_) );
OAI21X1 OAI21X1_667 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf5), .B(_2100__bF_buf1), .C(regs_5__1_), .Y(_2200_) );
OAI21X1 OAI21X1_668 ( .gnd(gnd), .vdd(vdd), .A(_1003__bF_buf2), .B(_2198__bF_buf3), .C(_2200_), .Y(_843_) );
OAI21X1 OAI21X1_669 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf4), .B(_2100__bF_buf0), .C(regs_5__2_), .Y(_2201_) );
OAI21X1 OAI21X1_670 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf2), .B(_2198__bF_buf2), .C(_2201_), .Y(_854_) );
OAI21X1 OAI21X1_671 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf3), .B(_2100__bF_buf8), .C(regs_5__3_), .Y(_2202_) );
OAI21X1 OAI21X1_672 ( .gnd(gnd), .vdd(vdd), .A(_1007__bF_buf2), .B(_2198__bF_buf1), .C(_2202_), .Y(_857_) );
OAI21X1 OAI21X1_673 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf2), .B(_2100__bF_buf7), .C(regs_5__4_), .Y(_2203_) );
OAI21X1 OAI21X1_674 ( .gnd(gnd), .vdd(vdd), .A(_1009__bF_buf1), .B(_2198__bF_buf0), .C(_2203_), .Y(_858_) );
OAI21X1 OAI21X1_675 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf1), .B(_2100__bF_buf6), .C(regs_5__5_), .Y(_2204_) );
OAI21X1 OAI21X1_676 ( .gnd(gnd), .vdd(vdd), .A(_1011__bF_buf1), .B(_2198__bF_buf4), .C(_2204_), .Y(_859_) );
OAI21X1 OAI21X1_677 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf0), .B(_2100__bF_buf5), .C(regs_5__6_), .Y(_2205_) );
OAI21X1 OAI21X1_678 ( .gnd(gnd), .vdd(vdd), .A(_1013__bF_buf1), .B(_2198__bF_buf3), .C(_2205_), .Y(_860_) );
OAI21X1 OAI21X1_679 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf10), .B(_2100__bF_buf4), .C(regs_5__7_), .Y(_2206_) );
OAI21X1 OAI21X1_680 ( .gnd(gnd), .vdd(vdd), .A(_1015__bF_buf1), .B(_2198__bF_buf2), .C(_2206_), .Y(_861_) );
OAI21X1 OAI21X1_681 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf9), .B(_2100__bF_buf3), .C(regs_5__8_), .Y(_2207_) );
OAI21X1 OAI21X1_682 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf1), .B(_2198__bF_buf1), .C(_2207_), .Y(_862_) );
OAI21X1 OAI21X1_683 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf8), .B(_2100__bF_buf2), .C(regs_5__9_), .Y(_2208_) );
OAI21X1 OAI21X1_684 ( .gnd(gnd), .vdd(vdd), .A(_1019__bF_buf1), .B(_2198__bF_buf0), .C(_2208_), .Y(_863_) );
OAI21X1 OAI21X1_685 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf7), .B(_2100__bF_buf1), .C(regs_5__10_), .Y(_2209_) );
OAI21X1 OAI21X1_686 ( .gnd(gnd), .vdd(vdd), .A(_1021__bF_buf1), .B(_2198__bF_buf4), .C(_2209_), .Y(_833_) );
OAI21X1 OAI21X1_687 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf6), .B(_2100__bF_buf0), .C(regs_5__11_), .Y(_2210_) );
OAI21X1 OAI21X1_688 ( .gnd(gnd), .vdd(vdd), .A(_1023__bF_buf1), .B(_2198__bF_buf3), .C(_2210_), .Y(_834_) );
OAI21X1 OAI21X1_689 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf5), .B(_2100__bF_buf8), .C(regs_5__12_), .Y(_2211_) );
OAI21X1 OAI21X1_690 ( .gnd(gnd), .vdd(vdd), .A(_1025__bF_buf1), .B(_2198__bF_buf2), .C(_2211_), .Y(_835_) );
OAI21X1 OAI21X1_691 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf4), .B(_2100__bF_buf7), .C(regs_5__13_), .Y(_2212_) );
OAI21X1 OAI21X1_692 ( .gnd(gnd), .vdd(vdd), .A(_1027__bF_buf1), .B(_2198__bF_buf1), .C(_2212_), .Y(_836_) );
OAI21X1 OAI21X1_693 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf3), .B(_2100__bF_buf6), .C(regs_5__14_), .Y(_2213_) );
OAI21X1 OAI21X1_694 ( .gnd(gnd), .vdd(vdd), .A(_1029__bF_buf1), .B(_2198__bF_buf0), .C(_2213_), .Y(_837_) );
OAI21X1 OAI21X1_695 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf2), .B(_2100__bF_buf5), .C(regs_5__15_), .Y(_2214_) );
OAI21X1 OAI21X1_696 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf1), .B(_2198__bF_buf4), .C(_2214_), .Y(_838_) );
OAI21X1 OAI21X1_697 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf1), .B(_2100__bF_buf4), .C(regs_5__16_), .Y(_2215_) );
OAI21X1 OAI21X1_698 ( .gnd(gnd), .vdd(vdd), .A(_1033__bF_buf1), .B(_2198__bF_buf3), .C(_2215_), .Y(_839_) );
OAI21X1 OAI21X1_699 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf0), .B(_2100__bF_buf3), .C(regs_5__17_), .Y(_2216_) );
OAI21X1 OAI21X1_700 ( .gnd(gnd), .vdd(vdd), .A(_1035__bF_buf1), .B(_2198__bF_buf2), .C(_2216_), .Y(_840_) );
OAI21X1 OAI21X1_701 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf10), .B(_2100__bF_buf2), .C(regs_5__18_), .Y(_2217_) );
OAI21X1 OAI21X1_702 ( .gnd(gnd), .vdd(vdd), .A(_1037__bF_buf1), .B(_2198__bF_buf1), .C(_2217_), .Y(_841_) );
OAI21X1 OAI21X1_703 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf9), .B(_2100__bF_buf1), .C(regs_5__19_), .Y(_2218_) );
OAI21X1 OAI21X1_704 ( .gnd(gnd), .vdd(vdd), .A(_1039__bF_buf1), .B(_2198__bF_buf0), .C(_2218_), .Y(_842_) );
OAI21X1 OAI21X1_705 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf8), .B(_2100__bF_buf0), .C(regs_5__20_), .Y(_2219_) );
OAI21X1 OAI21X1_706 ( .gnd(gnd), .vdd(vdd), .A(_1041__bF_buf1), .B(_2198__bF_buf4), .C(_2219_), .Y(_844_) );
OAI21X1 OAI21X1_707 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf7), .B(_2100__bF_buf8), .C(regs_5__21_), .Y(_2220_) );
OAI21X1 OAI21X1_708 ( .gnd(gnd), .vdd(vdd), .A(_1043__bF_buf1), .B(_2198__bF_buf3), .C(_2220_), .Y(_845_) );
OAI21X1 OAI21X1_709 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf6), .B(_2100__bF_buf7), .C(regs_5__22_), .Y(_2221_) );
OAI21X1 OAI21X1_710 ( .gnd(gnd), .vdd(vdd), .A(_1045__bF_buf1), .B(_2198__bF_buf2), .C(_2221_), .Y(_846_) );
OAI21X1 OAI21X1_711 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf5), .B(_2100__bF_buf6), .C(regs_5__23_), .Y(_2222_) );
OAI21X1 OAI21X1_712 ( .gnd(gnd), .vdd(vdd), .A(_1047__bF_buf1), .B(_2198__bF_buf1), .C(_2222_), .Y(_847_) );
OAI21X1 OAI21X1_713 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf4), .B(_2100__bF_buf5), .C(regs_5__24_), .Y(_2223_) );
OAI21X1 OAI21X1_714 ( .gnd(gnd), .vdd(vdd), .A(_1049__bF_buf1), .B(_2198__bF_buf0), .C(_2223_), .Y(_848_) );
OAI21X1 OAI21X1_715 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf3), .B(_2100__bF_buf4), .C(regs_5__25_), .Y(_2224_) );
OAI21X1 OAI21X1_716 ( .gnd(gnd), .vdd(vdd), .A(_1051__bF_buf1), .B(_2198__bF_buf4), .C(_2224_), .Y(_849_) );
OAI21X1 OAI21X1_717 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf2), .B(_2100__bF_buf3), .C(regs_5__26_), .Y(_2225_) );
OAI21X1 OAI21X1_718 ( .gnd(gnd), .vdd(vdd), .A(_1053__bF_buf1), .B(_2198__bF_buf3), .C(_2225_), .Y(_850_) );
OAI21X1 OAI21X1_719 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf1), .B(_2100__bF_buf2), .C(regs_5__27_), .Y(_2226_) );
OAI21X1 OAI21X1_720 ( .gnd(gnd), .vdd(vdd), .A(_1055__bF_buf1), .B(_2198__bF_buf2), .C(_2226_), .Y(_851_) );
OAI21X1 OAI21X1_721 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf0), .B(_2100__bF_buf1), .C(regs_5__28_), .Y(_2227_) );
OAI21X1 OAI21X1_722 ( .gnd(gnd), .vdd(vdd), .A(_1057__bF_buf1), .B(_2198__bF_buf1), .C(_2227_), .Y(_852_) );
OAI21X1 OAI21X1_723 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf10), .B(_2100__bF_buf0), .C(regs_5__29_), .Y(_2228_) );
OAI21X1 OAI21X1_724 ( .gnd(gnd), .vdd(vdd), .A(_1059__bF_buf1), .B(_2198__bF_buf0), .C(_2228_), .Y(_853_) );
OAI21X1 OAI21X1_725 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf9), .B(_2100__bF_buf8), .C(regs_5__30_), .Y(_2229_) );
OAI21X1 OAI21X1_726 ( .gnd(gnd), .vdd(vdd), .A(_1061__bF_buf1), .B(_2198__bF_buf4), .C(_2229_), .Y(_855_) );
OAI21X1 OAI21X1_727 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf8), .B(_2100__bF_buf7), .C(regs_5__31_), .Y(_2230_) );
OAI21X1 OAI21X1_728 ( .gnd(gnd), .vdd(vdd), .A(_1063__bF_buf1), .B(_2198__bF_buf3), .C(_2230_), .Y(_856_) );
NAND2X1 NAND2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_2099_), .B(_1273_), .Y(_2231_) );
OAI21X1 OAI21X1_729 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf6), .B(_1104__bF_buf4), .C(regs_4__0_), .Y(_2232_) );
OAI21X1 OAI21X1_730 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf4), .B(_992__bF_buf1), .C(_2232_), .Y(_800_) );
OAI21X1 OAI21X1_731 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf5), .B(_1104__bF_buf3), .C(regs_4__1_), .Y(_2233_) );
OAI21X1 OAI21X1_732 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf3), .B(_1003__bF_buf1), .C(_2233_), .Y(_811_) );
OAI21X1 OAI21X1_733 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf4), .B(_1104__bF_buf2), .C(regs_4__2_), .Y(_2234_) );
OAI21X1 OAI21X1_734 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf2), .B(_1005__bF_buf1), .C(_2234_), .Y(_822_) );
OAI21X1 OAI21X1_735 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf3), .B(_1104__bF_buf1), .C(regs_4__3_), .Y(_2235_) );
OAI21X1 OAI21X1_736 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf1), .B(_1007__bF_buf1), .C(_2235_), .Y(_825_) );
OAI21X1 OAI21X1_737 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf2), .B(_1104__bF_buf0), .C(regs_4__4_), .Y(_2236_) );
OAI21X1 OAI21X1_738 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf0), .B(_1009__bF_buf0), .C(_2236_), .Y(_826_) );
OAI21X1 OAI21X1_739 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf1), .B(_1104__bF_buf14), .C(regs_4__5_), .Y(_2237_) );
OAI21X1 OAI21X1_740 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf4), .B(_1011__bF_buf0), .C(_2237_), .Y(_827_) );
OAI21X1 OAI21X1_741 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf0), .B(_1104__bF_buf13), .C(regs_4__6_), .Y(_2238_) );
OAI21X1 OAI21X1_742 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf3), .B(_1013__bF_buf0), .C(_2238_), .Y(_828_) );
OAI21X1 OAI21X1_743 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf8), .B(_1104__bF_buf12), .C(regs_4__7_), .Y(_2239_) );
OAI21X1 OAI21X1_744 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf2), .B(_1015__bF_buf0), .C(_2239_), .Y(_829_) );
OAI21X1 OAI21X1_745 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf7), .B(_1104__bF_buf11), .C(regs_4__8_), .Y(_2240_) );
OAI21X1 OAI21X1_746 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf1), .B(_1017__bF_buf0), .C(_2240_), .Y(_830_) );
OAI21X1 OAI21X1_747 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf6), .B(_1104__bF_buf10), .C(regs_4__9_), .Y(_2241_) );
OAI21X1 OAI21X1_748 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf0), .B(_1019__bF_buf0), .C(_2241_), .Y(_831_) );
OAI21X1 OAI21X1_749 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf5), .B(_1104__bF_buf9), .C(regs_4__10_), .Y(_2242_) );
OAI21X1 OAI21X1_750 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf4), .B(_1021__bF_buf0), .C(_2242_), .Y(_801_) );
OAI21X1 OAI21X1_751 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf4), .B(_1104__bF_buf8), .C(regs_4__11_), .Y(_2243_) );
OAI21X1 OAI21X1_752 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf3), .B(_1023__bF_buf0), .C(_2243_), .Y(_802_) );
OAI21X1 OAI21X1_753 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf3), .B(_1104__bF_buf7), .C(regs_4__12_), .Y(_2244_) );
OAI21X1 OAI21X1_754 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf2), .B(_1025__bF_buf0), .C(_2244_), .Y(_803_) );
OAI21X1 OAI21X1_755 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf2), .B(_1104__bF_buf6), .C(regs_4__13_), .Y(_2245_) );
OAI21X1 OAI21X1_756 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf1), .B(_1027__bF_buf0), .C(_2245_), .Y(_804_) );
OAI21X1 OAI21X1_757 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf1), .B(_1104__bF_buf5), .C(regs_4__14_), .Y(_2246_) );
OAI21X1 OAI21X1_758 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf0), .B(_1029__bF_buf0), .C(_2246_), .Y(_805_) );
OAI21X1 OAI21X1_759 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf0), .B(_1104__bF_buf4), .C(regs_4__15_), .Y(_2247_) );
OAI21X1 OAI21X1_760 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf4), .B(_1031__bF_buf0), .C(_2247_), .Y(_806_) );
OAI21X1 OAI21X1_761 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf8), .B(_1104__bF_buf3), .C(regs_4__16_), .Y(_2248_) );
OAI21X1 OAI21X1_762 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf3), .B(_1033__bF_buf0), .C(_2248_), .Y(_807_) );
OAI21X1 OAI21X1_763 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf7), .B(_1104__bF_buf2), .C(regs_4__17_), .Y(_2249_) );
OAI21X1 OAI21X1_764 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf2), .B(_1035__bF_buf0), .C(_2249_), .Y(_808_) );
OAI21X1 OAI21X1_765 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf6), .B(_1104__bF_buf1), .C(regs_4__18_), .Y(_2250_) );
OAI21X1 OAI21X1_766 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf1), .B(_1037__bF_buf0), .C(_2250_), .Y(_809_) );
OAI21X1 OAI21X1_767 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf5), .B(_1104__bF_buf0), .C(regs_4__19_), .Y(_2251_) );
OAI21X1 OAI21X1_768 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf0), .B(_1039__bF_buf0), .C(_2251_), .Y(_810_) );
OAI21X1 OAI21X1_769 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf4), .B(_1104__bF_buf14), .C(regs_4__20_), .Y(_2252_) );
OAI21X1 OAI21X1_770 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf4), .B(_1041__bF_buf0), .C(_2252_), .Y(_812_) );
OAI21X1 OAI21X1_771 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf3), .B(_1104__bF_buf13), .C(regs_4__21_), .Y(_2253_) );
OAI21X1 OAI21X1_772 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf3), .B(_1043__bF_buf0), .C(_2253_), .Y(_813_) );
OAI21X1 OAI21X1_773 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf2), .B(_1104__bF_buf12), .C(regs_4__22_), .Y(_2254_) );
OAI21X1 OAI21X1_774 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf2), .B(_1045__bF_buf0), .C(_2254_), .Y(_814_) );
OAI21X1 OAI21X1_775 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf1), .B(_1104__bF_buf11), .C(regs_4__23_), .Y(_2255_) );
OAI21X1 OAI21X1_776 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf1), .B(_1047__bF_buf0), .C(_2255_), .Y(_815_) );
OAI21X1 OAI21X1_777 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf0), .B(_1104__bF_buf10), .C(regs_4__24_), .Y(_2256_) );
OAI21X1 OAI21X1_778 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf0), .B(_1049__bF_buf0), .C(_2256_), .Y(_816_) );
OAI21X1 OAI21X1_779 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf8), .B(_1104__bF_buf9), .C(regs_4__25_), .Y(_2257_) );
OAI21X1 OAI21X1_780 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf4), .B(_1051__bF_buf0), .C(_2257_), .Y(_817_) );
OAI21X1 OAI21X1_781 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf7), .B(_1104__bF_buf8), .C(regs_4__26_), .Y(_2258_) );
OAI21X1 OAI21X1_782 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf3), .B(_1053__bF_buf0), .C(_2258_), .Y(_818_) );
OAI21X1 OAI21X1_783 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf6), .B(_1104__bF_buf7), .C(regs_4__27_), .Y(_2259_) );
OAI21X1 OAI21X1_784 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf2), .B(_1055__bF_buf0), .C(_2259_), .Y(_819_) );
OAI21X1 OAI21X1_785 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf5), .B(_1104__bF_buf6), .C(regs_4__28_), .Y(_2260_) );
OAI21X1 OAI21X1_786 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf1), .B(_1057__bF_buf0), .C(_2260_), .Y(_820_) );
OAI21X1 OAI21X1_787 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf4), .B(_1104__bF_buf5), .C(regs_4__29_), .Y(_2261_) );
OAI21X1 OAI21X1_788 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf0), .B(_1059__bF_buf0), .C(_2261_), .Y(_821_) );
OAI21X1 OAI21X1_789 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf3), .B(_1104__bF_buf4), .C(regs_4__30_), .Y(_2262_) );
OAI21X1 OAI21X1_790 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf4), .B(_1061__bF_buf0), .C(_2262_), .Y(_823_) );
OAI21X1 OAI21X1_791 ( .gnd(gnd), .vdd(vdd), .A(_2100__bF_buf2), .B(_1104__bF_buf3), .C(regs_4__31_), .Y(_2263_) );
OAI21X1 OAI21X1_792 ( .gnd(gnd), .vdd(vdd), .A(_2231__bF_buf3), .B(_1063__bF_buf0), .C(_2263_), .Y(_824_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_2098_), .B(_1139_), .Y(_2264_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf10), .B(_1142__bF_buf0), .Y(_2265_) );
OAI21X1 OAI21X1_793 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf9), .B(_1142__bF_buf5), .C(regs_3__0_), .Y(_2266_) );
OAI21X1 OAI21X1_794 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf4), .B(_992__bF_buf0), .C(_2266_), .Y(_768_) );
OAI21X1 OAI21X1_795 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf8), .B(_1142__bF_buf4), .C(regs_3__1_), .Y(_2267_) );
OAI21X1 OAI21X1_796 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf3), .B(_1003__bF_buf0), .C(_2267_), .Y(_779_) );
OAI21X1 OAI21X1_797 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf7), .B(_1142__bF_buf3), .C(regs_3__2_), .Y(_2268_) );
OAI21X1 OAI21X1_798 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf2), .B(_1005__bF_buf0), .C(_2268_), .Y(_790_) );
OAI21X1 OAI21X1_799 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf6), .B(_1142__bF_buf2), .C(regs_3__3_), .Y(_2269_) );
OAI21X1 OAI21X1_800 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf1), .B(_1007__bF_buf0), .C(_2269_), .Y(_793_) );
OAI21X1 OAI21X1_801 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf5), .B(_1142__bF_buf1), .C(regs_3__4_), .Y(_2270_) );
OAI21X1 OAI21X1_802 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf0), .B(_1009__bF_buf3), .C(_2270_), .Y(_794_) );
OAI21X1 OAI21X1_803 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf4), .B(_1142__bF_buf0), .C(regs_3__5_), .Y(_2271_) );
OAI21X1 OAI21X1_804 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf4), .B(_1011__bF_buf3), .C(_2271_), .Y(_795_) );
OAI21X1 OAI21X1_805 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf3), .B(_1142__bF_buf5), .C(regs_3__6_), .Y(_2272_) );
OAI21X1 OAI21X1_806 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf3), .B(_1013__bF_buf3), .C(_2272_), .Y(_796_) );
OAI21X1 OAI21X1_807 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf2), .B(_1142__bF_buf4), .C(regs_3__7_), .Y(_2273_) );
OAI21X1 OAI21X1_808 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf2), .B(_1015__bF_buf3), .C(_2273_), .Y(_797_) );
OAI21X1 OAI21X1_809 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf1), .B(_1142__bF_buf3), .C(regs_3__8_), .Y(_2274_) );
OAI21X1 OAI21X1_810 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf1), .B(_1017__bF_buf3), .C(_2274_), .Y(_798_) );
OAI21X1 OAI21X1_811 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf0), .B(_1142__bF_buf2), .C(regs_3__9_), .Y(_2275_) );
OAI21X1 OAI21X1_812 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf0), .B(_1019__bF_buf3), .C(_2275_), .Y(_799_) );
OAI21X1 OAI21X1_813 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf10), .B(_1142__bF_buf1), .C(regs_3__10_), .Y(_2276_) );
OAI21X1 OAI21X1_814 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf4), .B(_1021__bF_buf3), .C(_2276_), .Y(_769_) );
OAI21X1 OAI21X1_815 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf9), .B(_1142__bF_buf0), .C(regs_3__11_), .Y(_2277_) );
OAI21X1 OAI21X1_816 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf3), .B(_1023__bF_buf3), .C(_2277_), .Y(_770_) );
OAI21X1 OAI21X1_817 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf8), .B(_1142__bF_buf5), .C(regs_3__12_), .Y(_2278_) );
OAI21X1 OAI21X1_818 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf2), .B(_1025__bF_buf3), .C(_2278_), .Y(_771_) );
OAI21X1 OAI21X1_819 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf7), .B(_1142__bF_buf4), .C(regs_3__13_), .Y(_2279_) );
OAI21X1 OAI21X1_820 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf1), .B(_1027__bF_buf3), .C(_2279_), .Y(_772_) );
OAI21X1 OAI21X1_821 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf6), .B(_1142__bF_buf3), .C(regs_3__14_), .Y(_2280_) );
OAI21X1 OAI21X1_822 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf0), .B(_1029__bF_buf3), .C(_2280_), .Y(_773_) );
OAI21X1 OAI21X1_823 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf5), .B(_1142__bF_buf2), .C(regs_3__15_), .Y(_2281_) );
OAI21X1 OAI21X1_824 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf4), .B(_1031__bF_buf3), .C(_2281_), .Y(_774_) );
OAI21X1 OAI21X1_825 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf4), .B(_1142__bF_buf1), .C(regs_3__16_), .Y(_2282_) );
OAI21X1 OAI21X1_826 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf3), .B(_1033__bF_buf3), .C(_2282_), .Y(_775_) );
OAI21X1 OAI21X1_827 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf3), .B(_1142__bF_buf0), .C(regs_3__17_), .Y(_2283_) );
OAI21X1 OAI21X1_828 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf2), .B(_1035__bF_buf3), .C(_2283_), .Y(_776_) );
OAI21X1 OAI21X1_829 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf2), .B(_1142__bF_buf5), .C(regs_3__18_), .Y(_2284_) );
OAI21X1 OAI21X1_830 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf1), .B(_1037__bF_buf3), .C(_2284_), .Y(_777_) );
OAI21X1 OAI21X1_831 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf1), .B(_1142__bF_buf4), .C(regs_3__19_), .Y(_2285_) );
OAI21X1 OAI21X1_832 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf0), .B(_1039__bF_buf3), .C(_2285_), .Y(_778_) );
OAI21X1 OAI21X1_833 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf0), .B(_1142__bF_buf3), .C(regs_3__20_), .Y(_2286_) );
OAI21X1 OAI21X1_834 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf4), .B(_1041__bF_buf3), .C(_2286_), .Y(_780_) );
OAI21X1 OAI21X1_835 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf10), .B(_1142__bF_buf2), .C(regs_3__21_), .Y(_2287_) );
OAI21X1 OAI21X1_836 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf3), .B(_1043__bF_buf3), .C(_2287_), .Y(_781_) );
OAI21X1 OAI21X1_837 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf9), .B(_1142__bF_buf1), .C(regs_3__22_), .Y(_2288_) );
OAI21X1 OAI21X1_838 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf2), .B(_1045__bF_buf3), .C(_2288_), .Y(_782_) );
OAI21X1 OAI21X1_839 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf8), .B(_1142__bF_buf0), .C(regs_3__23_), .Y(_2289_) );
OAI21X1 OAI21X1_840 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf1), .B(_1047__bF_buf3), .C(_2289_), .Y(_783_) );
OAI21X1 OAI21X1_841 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf7), .B(_1142__bF_buf5), .C(regs_3__24_), .Y(_2290_) );
OAI21X1 OAI21X1_842 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf0), .B(_1049__bF_buf3), .C(_2290_), .Y(_784_) );
OAI21X1 OAI21X1_843 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf6), .B(_1142__bF_buf4), .C(regs_3__25_), .Y(_2291_) );
OAI21X1 OAI21X1_844 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf4), .B(_1051__bF_buf3), .C(_2291_), .Y(_785_) );
OAI21X1 OAI21X1_845 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf5), .B(_1142__bF_buf3), .C(regs_3__26_), .Y(_2292_) );
OAI21X1 OAI21X1_846 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf3), .B(_1053__bF_buf3), .C(_2292_), .Y(_786_) );
OAI21X1 OAI21X1_847 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf4), .B(_1142__bF_buf2), .C(regs_3__27_), .Y(_2293_) );
OAI21X1 OAI21X1_848 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf2), .B(_1055__bF_buf3), .C(_2293_), .Y(_787_) );
OAI21X1 OAI21X1_849 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf3), .B(_1142__bF_buf1), .C(regs_3__28_), .Y(_2294_) );
OAI21X1 OAI21X1_850 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf1), .B(_1057__bF_buf3), .C(_2294_), .Y(_788_) );
OAI21X1 OAI21X1_851 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf2), .B(_1142__bF_buf0), .C(regs_3__29_), .Y(_2295_) );
OAI21X1 OAI21X1_852 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf0), .B(_1059__bF_buf3), .C(_2295_), .Y(_789_) );
OAI21X1 OAI21X1_853 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf1), .B(_1142__bF_buf5), .C(regs_3__30_), .Y(_2296_) );
OAI21X1 OAI21X1_854 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf4), .B(_1061__bF_buf3), .C(_2296_), .Y(_791_) );
OAI21X1 OAI21X1_855 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf0), .B(_1142__bF_buf4), .C(regs_3__31_), .Y(_2297_) );
OAI21X1 OAI21X1_856 ( .gnd(gnd), .vdd(vdd), .A(_2265__bF_buf3), .B(_1063__bF_buf3), .C(_2297_), .Y(_792_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_2264__bF_buf10), .Y(_2298_) );
NAND2X1 NAND2X1_295 ( .gnd(gnd), .vdd(vdd), .A(_998_), .B(_2298_), .Y(_2299_) );
OAI21X1 OAI21X1_857 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf3), .B(_2264__bF_buf9), .C(regs_2__0_), .Y(_2300_) );
OAI21X1 OAI21X1_858 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf4), .B(_992__bF_buf3), .C(_2300_), .Y(_704_) );
OAI21X1 OAI21X1_859 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf2), .B(_2264__bF_buf8), .C(regs_2__1_), .Y(_2301_) );
OAI21X1 OAI21X1_860 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf3), .B(_1003__bF_buf3), .C(_2301_), .Y(_715_) );
OAI21X1 OAI21X1_861 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf1), .B(_2264__bF_buf7), .C(regs_2__2_), .Y(_2302_) );
OAI21X1 OAI21X1_862 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf2), .B(_1005__bF_buf3), .C(_2302_), .Y(_726_) );
OAI21X1 OAI21X1_863 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf0), .B(_2264__bF_buf6), .C(regs_2__3_), .Y(_2303_) );
OAI21X1 OAI21X1_864 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf1), .B(_1007__bF_buf3), .C(_2303_), .Y(_729_) );
OAI21X1 OAI21X1_865 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf9), .B(_2264__bF_buf5), .C(regs_2__4_), .Y(_2304_) );
OAI21X1 OAI21X1_866 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf0), .B(_1009__bF_buf2), .C(_2304_), .Y(_730_) );
OAI21X1 OAI21X1_867 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf8), .B(_2264__bF_buf4), .C(regs_2__5_), .Y(_2305_) );
OAI21X1 OAI21X1_868 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf4), .B(_1011__bF_buf2), .C(_2305_), .Y(_731_) );
OAI21X1 OAI21X1_869 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf7), .B(_2264__bF_buf3), .C(regs_2__6_), .Y(_2306_) );
OAI21X1 OAI21X1_870 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf3), .B(_1013__bF_buf2), .C(_2306_), .Y(_732_) );
OAI21X1 OAI21X1_871 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf6), .B(_2264__bF_buf2), .C(regs_2__7_), .Y(_2307_) );
OAI21X1 OAI21X1_872 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf2), .B(_1015__bF_buf2), .C(_2307_), .Y(_733_) );
OAI21X1 OAI21X1_873 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf5), .B(_2264__bF_buf1), .C(regs_2__8_), .Y(_2308_) );
OAI21X1 OAI21X1_874 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf1), .B(_1017__bF_buf2), .C(_2308_), .Y(_734_) );
OAI21X1 OAI21X1_875 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf4), .B(_2264__bF_buf0), .C(regs_2__9_), .Y(_2309_) );
OAI21X1 OAI21X1_876 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf0), .B(_1019__bF_buf2), .C(_2309_), .Y(_735_) );
OAI21X1 OAI21X1_877 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf3), .B(_2264__bF_buf10), .C(regs_2__10_), .Y(_2310_) );
OAI21X1 OAI21X1_878 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf4), .B(_1021__bF_buf2), .C(_2310_), .Y(_705_) );
OAI21X1 OAI21X1_879 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf2), .B(_2264__bF_buf9), .C(regs_2__11_), .Y(_2311_) );
OAI21X1 OAI21X1_880 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf3), .B(_1023__bF_buf2), .C(_2311_), .Y(_706_) );
OAI21X1 OAI21X1_881 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf1), .B(_2264__bF_buf8), .C(regs_2__12_), .Y(_2312_) );
OAI21X1 OAI21X1_882 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf2), .B(_1025__bF_buf2), .C(_2312_), .Y(_707_) );
OAI21X1 OAI21X1_883 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf0), .B(_2264__bF_buf7), .C(regs_2__13_), .Y(_2313_) );
OAI21X1 OAI21X1_884 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf1), .B(_1027__bF_buf2), .C(_2313_), .Y(_708_) );
OAI21X1 OAI21X1_885 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf9), .B(_2264__bF_buf6), .C(regs_2__14_), .Y(_2314_) );
OAI21X1 OAI21X1_886 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf0), .B(_1029__bF_buf2), .C(_2314_), .Y(_709_) );
OAI21X1 OAI21X1_887 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf8), .B(_2264__bF_buf5), .C(regs_2__15_), .Y(_2315_) );
OAI21X1 OAI21X1_888 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf4), .B(_1031__bF_buf2), .C(_2315_), .Y(_710_) );
OAI21X1 OAI21X1_889 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf7), .B(_2264__bF_buf4), .C(regs_2__16_), .Y(_2316_) );
OAI21X1 OAI21X1_890 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf3), .B(_1033__bF_buf2), .C(_2316_), .Y(_711_) );
OAI21X1 OAI21X1_891 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf6), .B(_2264__bF_buf3), .C(regs_2__17_), .Y(_2317_) );
OAI21X1 OAI21X1_892 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf2), .B(_1035__bF_buf2), .C(_2317_), .Y(_712_) );
OAI21X1 OAI21X1_893 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf5), .B(_2264__bF_buf2), .C(regs_2__18_), .Y(_2318_) );
OAI21X1 OAI21X1_894 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf1), .B(_1037__bF_buf2), .C(_2318_), .Y(_713_) );
OAI21X1 OAI21X1_895 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf4), .B(_2264__bF_buf1), .C(regs_2__19_), .Y(_2319_) );
OAI21X1 OAI21X1_896 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf0), .B(_1039__bF_buf2), .C(_2319_), .Y(_714_) );
OAI21X1 OAI21X1_897 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf3), .B(_2264__bF_buf0), .C(regs_2__20_), .Y(_2320_) );
OAI21X1 OAI21X1_898 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf4), .B(_1041__bF_buf2), .C(_2320_), .Y(_716_) );
OAI21X1 OAI21X1_899 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf2), .B(_2264__bF_buf10), .C(regs_2__21_), .Y(_2321_) );
OAI21X1 OAI21X1_900 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf3), .B(_1043__bF_buf2), .C(_2321_), .Y(_717_) );
OAI21X1 OAI21X1_901 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf1), .B(_2264__bF_buf9), .C(regs_2__22_), .Y(_2322_) );
OAI21X1 OAI21X1_902 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf2), .B(_1045__bF_buf2), .C(_2322_), .Y(_718_) );
OAI21X1 OAI21X1_903 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf0), .B(_2264__bF_buf8), .C(regs_2__23_), .Y(_2323_) );
OAI21X1 OAI21X1_904 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf1), .B(_1047__bF_buf2), .C(_2323_), .Y(_719_) );
OAI21X1 OAI21X1_905 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf9), .B(_2264__bF_buf7), .C(regs_2__24_), .Y(_2324_) );
OAI21X1 OAI21X1_906 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf0), .B(_1049__bF_buf2), .C(_2324_), .Y(_720_) );
OAI21X1 OAI21X1_907 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf8), .B(_2264__bF_buf6), .C(regs_2__25_), .Y(_2325_) );
OAI21X1 OAI21X1_908 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf4), .B(_1051__bF_buf2), .C(_2325_), .Y(_721_) );
OAI21X1 OAI21X1_909 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf7), .B(_2264__bF_buf5), .C(regs_2__26_), .Y(_2326_) );
OAI21X1 OAI21X1_910 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf3), .B(_1053__bF_buf2), .C(_2326_), .Y(_722_) );
OAI21X1 OAI21X1_911 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf6), .B(_2264__bF_buf4), .C(regs_2__27_), .Y(_2327_) );
OAI21X1 OAI21X1_912 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf2), .B(_1055__bF_buf2), .C(_2327_), .Y(_723_) );
OAI21X1 OAI21X1_913 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf5), .B(_2264__bF_buf3), .C(regs_2__28_), .Y(_2328_) );
OAI21X1 OAI21X1_914 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf1), .B(_1057__bF_buf2), .C(_2328_), .Y(_724_) );
OAI21X1 OAI21X1_915 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf4), .B(_2264__bF_buf2), .C(regs_2__29_), .Y(_2329_) );
OAI21X1 OAI21X1_916 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf0), .B(_1059__bF_buf2), .C(_2329_), .Y(_725_) );
OAI21X1 OAI21X1_917 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf3), .B(_2264__bF_buf1), .C(regs_2__30_), .Y(_2330_) );
OAI21X1 OAI21X1_918 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf4), .B(_1061__bF_buf2), .C(_2330_), .Y(_727_) );
OAI21X1 OAI21X1_919 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf2), .B(_2264__bF_buf0), .C(regs_2__31_), .Y(_2331_) );
OAI21X1 OAI21X1_920 ( .gnd(gnd), .vdd(vdd), .A(_2299__bF_buf3), .B(_1063__bF_buf2), .C(_2331_), .Y(_728_) );
NAND2X1 NAND2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_2298_), .Y(_2332_) );
OAI21X1 OAI21X1_921 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf7), .B(_2264__bF_buf10), .C(regs_1__0_), .Y(_2333_) );
OAI21X1 OAI21X1_922 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf4), .B(_992__bF_buf2), .C(_2333_), .Y(_352_) );
OAI21X1 OAI21X1_923 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf6), .B(_2264__bF_buf9), .C(regs_1__1_), .Y(_2334_) );
OAI21X1 OAI21X1_924 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf3), .B(_1003__bF_buf2), .C(_2334_), .Y(_363_) );
OAI21X1 OAI21X1_925 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf5), .B(_2264__bF_buf8), .C(regs_1__2_), .Y(_2335_) );
OAI21X1 OAI21X1_926 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf2), .B(_1005__bF_buf2), .C(_2335_), .Y(_374_) );
OAI21X1 OAI21X1_927 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf4), .B(_2264__bF_buf7), .C(regs_1__3_), .Y(_2336_) );
OAI21X1 OAI21X1_928 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf1), .B(_1007__bF_buf2), .C(_2336_), .Y(_377_) );
OAI21X1 OAI21X1_929 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf3), .B(_2264__bF_buf6), .C(regs_1__4_), .Y(_2337_) );
OAI21X1 OAI21X1_930 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf0), .B(_1009__bF_buf1), .C(_2337_), .Y(_378_) );
OAI21X1 OAI21X1_931 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf2), .B(_2264__bF_buf5), .C(regs_1__5_), .Y(_2338_) );
OAI21X1 OAI21X1_932 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf4), .B(_1011__bF_buf1), .C(_2338_), .Y(_379_) );
OAI21X1 OAI21X1_933 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf1), .B(_2264__bF_buf4), .C(regs_1__6_), .Y(_2339_) );
OAI21X1 OAI21X1_934 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf3), .B(_1013__bF_buf1), .C(_2339_), .Y(_380_) );
OAI21X1 OAI21X1_935 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf0), .B(_2264__bF_buf3), .C(regs_1__7_), .Y(_2340_) );
OAI21X1 OAI21X1_936 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf2), .B(_1015__bF_buf1), .C(_2340_), .Y(_381_) );
OAI21X1 OAI21X1_937 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf10), .B(_2264__bF_buf2), .C(regs_1__8_), .Y(_2341_) );
OAI21X1 OAI21X1_938 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf1), .B(_1017__bF_buf1), .C(_2341_), .Y(_382_) );
OAI21X1 OAI21X1_939 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf9), .B(_2264__bF_buf1), .C(regs_1__9_), .Y(_2342_) );
OAI21X1 OAI21X1_940 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf0), .B(_1019__bF_buf1), .C(_2342_), .Y(_383_) );
OAI21X1 OAI21X1_941 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf8), .B(_2264__bF_buf0), .C(regs_1__10_), .Y(_2343_) );
OAI21X1 OAI21X1_942 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf4), .B(_1021__bF_buf1), .C(_2343_), .Y(_353_) );
OAI21X1 OAI21X1_943 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf7), .B(_2264__bF_buf10), .C(regs_1__11_), .Y(_2344_) );
OAI21X1 OAI21X1_944 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf3), .B(_1023__bF_buf1), .C(_2344_), .Y(_354_) );
OAI21X1 OAI21X1_945 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf6), .B(_2264__bF_buf9), .C(regs_1__12_), .Y(_2345_) );
OAI21X1 OAI21X1_946 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf2), .B(_1025__bF_buf1), .C(_2345_), .Y(_355_) );
OAI21X1 OAI21X1_947 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf5), .B(_2264__bF_buf8), .C(regs_1__13_), .Y(_2346_) );
OAI21X1 OAI21X1_948 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf1), .B(_1027__bF_buf1), .C(_2346_), .Y(_356_) );
OAI21X1 OAI21X1_949 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf4), .B(_2264__bF_buf7), .C(regs_1__14_), .Y(_2347_) );
OAI21X1 OAI21X1_950 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf0), .B(_1029__bF_buf1), .C(_2347_), .Y(_357_) );
OAI21X1 OAI21X1_951 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf3), .B(_2264__bF_buf6), .C(regs_1__15_), .Y(_2348_) );
OAI21X1 OAI21X1_952 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf4), .B(_1031__bF_buf1), .C(_2348_), .Y(_358_) );
OAI21X1 OAI21X1_953 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf2), .B(_2264__bF_buf5), .C(regs_1__16_), .Y(_2349_) );
OAI21X1 OAI21X1_954 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf3), .B(_1033__bF_buf1), .C(_2349_), .Y(_359_) );
OAI21X1 OAI21X1_955 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf1), .B(_2264__bF_buf4), .C(regs_1__17_), .Y(_2350_) );
OAI21X1 OAI21X1_956 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf2), .B(_1035__bF_buf1), .C(_2350_), .Y(_360_) );
OAI21X1 OAI21X1_957 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf0), .B(_2264__bF_buf3), .C(regs_1__18_), .Y(_2351_) );
OAI21X1 OAI21X1_958 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf1), .B(_1037__bF_buf1), .C(_2351_), .Y(_361_) );
OAI21X1 OAI21X1_959 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf10), .B(_2264__bF_buf2), .C(regs_1__19_), .Y(_2352_) );
OAI21X1 OAI21X1_960 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf0), .B(_1039__bF_buf1), .C(_2352_), .Y(_362_) );
OAI21X1 OAI21X1_961 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf9), .B(_2264__bF_buf1), .C(regs_1__20_), .Y(_2353_) );
OAI21X1 OAI21X1_962 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf4), .B(_1041__bF_buf1), .C(_2353_), .Y(_364_) );
OAI21X1 OAI21X1_963 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf8), .B(_2264__bF_buf0), .C(regs_1__21_), .Y(_2354_) );
OAI21X1 OAI21X1_964 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf3), .B(_1043__bF_buf1), .C(_2354_), .Y(_365_) );
OAI21X1 OAI21X1_965 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf7), .B(_2264__bF_buf10), .C(regs_1__22_), .Y(_2355_) );
OAI21X1 OAI21X1_966 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf2), .B(_1045__bF_buf1), .C(_2355_), .Y(_366_) );
OAI21X1 OAI21X1_967 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf6), .B(_2264__bF_buf9), .C(regs_1__23_), .Y(_2356_) );
OAI21X1 OAI21X1_968 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf1), .B(_1047__bF_buf1), .C(_2356_), .Y(_367_) );
OAI21X1 OAI21X1_969 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf5), .B(_2264__bF_buf8), .C(regs_1__24_), .Y(_2357_) );
OAI21X1 OAI21X1_970 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf0), .B(_1049__bF_buf1), .C(_2357_), .Y(_368_) );
OAI21X1 OAI21X1_971 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf4), .B(_2264__bF_buf7), .C(regs_1__25_), .Y(_2358_) );
OAI21X1 OAI21X1_972 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf4), .B(_1051__bF_buf1), .C(_2358_), .Y(_369_) );
OAI21X1 OAI21X1_973 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf3), .B(_2264__bF_buf6), .C(regs_1__26_), .Y(_2359_) );
OAI21X1 OAI21X1_974 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf3), .B(_1053__bF_buf1), .C(_2359_), .Y(_370_) );
OAI21X1 OAI21X1_975 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf2), .B(_2264__bF_buf5), .C(regs_1__27_), .Y(_2360_) );
OAI21X1 OAI21X1_976 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf2), .B(_1055__bF_buf1), .C(_2360_), .Y(_371_) );
OAI21X1 OAI21X1_977 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf1), .B(_2264__bF_buf4), .C(regs_1__28_), .Y(_2361_) );
OAI21X1 OAI21X1_978 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf1), .B(_1057__bF_buf1), .C(_2361_), .Y(_372_) );
OAI21X1 OAI21X1_979 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf0), .B(_2264__bF_buf3), .C(regs_1__29_), .Y(_2362_) );
OAI21X1 OAI21X1_980 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf0), .B(_1059__bF_buf1), .C(_2362_), .Y(_373_) );
OAI21X1 OAI21X1_981 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf10), .B(_2264__bF_buf2), .C(regs_1__30_), .Y(_2363_) );
OAI21X1 OAI21X1_982 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf4), .B(_1061__bF_buf1), .C(_2363_), .Y(_375_) );
OAI21X1 OAI21X1_983 ( .gnd(gnd), .vdd(vdd), .A(_1070__bF_buf9), .B(_2264__bF_buf1), .C(regs_1__31_), .Y(_2364_) );
OAI21X1 OAI21X1_984 ( .gnd(gnd), .vdd(vdd), .A(_2332__bF_buf3), .B(_1063__bF_buf1), .C(_2364_), .Y(_376_) );
NAND2X1 NAND2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_1273_), .B(_2298_), .Y(_2365_) );
OAI21X1 OAI21X1_985 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf2), .B(_2264__bF_buf0), .C(regs_0__0_), .Y(_2366_) );
OAI21X1 OAI21X1_986 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf4), .B(_992__bF_buf1), .C(_2366_), .Y(_0_) );
OAI21X1 OAI21X1_987 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf1), .B(_2264__bF_buf10), .C(regs_0__1_), .Y(_2367_) );
OAI21X1 OAI21X1_988 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf3), .B(_1003__bF_buf1), .C(_2367_), .Y(_11_) );
OAI21X1 OAI21X1_989 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf0), .B(_2264__bF_buf9), .C(regs_0__2_), .Y(_2368_) );
OAI21X1 OAI21X1_990 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf2), .B(_1005__bF_buf1), .C(_2368_), .Y(_22_) );
OAI21X1 OAI21X1_991 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf14), .B(_2264__bF_buf8), .C(regs_0__3_), .Y(_2369_) );
OAI21X1 OAI21X1_992 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf1), .B(_1007__bF_buf1), .C(_2369_), .Y(_25_) );
OAI21X1 OAI21X1_993 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf13), .B(_2264__bF_buf7), .C(regs_0__4_), .Y(_2370_) );
OAI21X1 OAI21X1_994 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf0), .B(_1009__bF_buf0), .C(_2370_), .Y(_26_) );
OAI21X1 OAI21X1_995 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf12), .B(_2264__bF_buf6), .C(regs_0__5_), .Y(_2371_) );
OAI21X1 OAI21X1_996 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf4), .B(_1011__bF_buf0), .C(_2371_), .Y(_27_) );
OAI21X1 OAI21X1_997 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf11), .B(_2264__bF_buf5), .C(regs_0__6_), .Y(_2372_) );
OAI21X1 OAI21X1_998 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf3), .B(_1013__bF_buf0), .C(_2372_), .Y(_28_) );
OAI21X1 OAI21X1_999 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf10), .B(_2264__bF_buf4), .C(regs_0__7_), .Y(_2373_) );
OAI21X1 OAI21X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf2), .B(_1015__bF_buf0), .C(_2373_), .Y(_29_) );
OAI21X1 OAI21X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf9), .B(_2264__bF_buf3), .C(regs_0__8_), .Y(_2374_) );
OAI21X1 OAI21X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf1), .B(_1017__bF_buf0), .C(_2374_), .Y(_30_) );
OAI21X1 OAI21X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf8), .B(_2264__bF_buf2), .C(regs_0__9_), .Y(_2375_) );
OAI21X1 OAI21X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf0), .B(_1019__bF_buf0), .C(_2375_), .Y(_31_) );
OAI21X1 OAI21X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf7), .B(_2264__bF_buf1), .C(regs_0__10_), .Y(_2376_) );
OAI21X1 OAI21X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf4), .B(_1021__bF_buf0), .C(_2376_), .Y(_1_) );
OAI21X1 OAI21X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf6), .B(_2264__bF_buf0), .C(regs_0__11_), .Y(_2377_) );
OAI21X1 OAI21X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf3), .B(_1023__bF_buf0), .C(_2377_), .Y(_2_) );
OAI21X1 OAI21X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf5), .B(_2264__bF_buf10), .C(regs_0__12_), .Y(_2378_) );
OAI21X1 OAI21X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf2), .B(_1025__bF_buf0), .C(_2378_), .Y(_3_) );
OAI21X1 OAI21X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf4), .B(_2264__bF_buf9), .C(regs_0__13_), .Y(_2379_) );
OAI21X1 OAI21X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf1), .B(_1027__bF_buf0), .C(_2379_), .Y(_4_) );
OAI21X1 OAI21X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf3), .B(_2264__bF_buf8), .C(regs_0__14_), .Y(_2380_) );
OAI21X1 OAI21X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf0), .B(_1029__bF_buf0), .C(_2380_), .Y(_5_) );
OAI21X1 OAI21X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf2), .B(_2264__bF_buf7), .C(regs_0__15_), .Y(_2381_) );
OAI21X1 OAI21X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf4), .B(_1031__bF_buf0), .C(_2381_), .Y(_6_) );
OAI21X1 OAI21X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf1), .B(_2264__bF_buf6), .C(regs_0__16_), .Y(_2382_) );
OAI21X1 OAI21X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf3), .B(_1033__bF_buf0), .C(_2382_), .Y(_7_) );
OAI21X1 OAI21X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf0), .B(_2264__bF_buf5), .C(regs_0__17_), .Y(_2383_) );
OAI21X1 OAI21X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf2), .B(_1035__bF_buf0), .C(_2383_), .Y(_8_) );
OAI21X1 OAI21X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf14), .B(_2264__bF_buf4), .C(regs_0__18_), .Y(_2384_) );
OAI21X1 OAI21X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf1), .B(_1037__bF_buf0), .C(_2384_), .Y(_9_) );
OAI21X1 OAI21X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf13), .B(_2264__bF_buf3), .C(regs_0__19_), .Y(_2385_) );
OAI21X1 OAI21X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf0), .B(_1039__bF_buf0), .C(_2385_), .Y(_10_) );
OAI21X1 OAI21X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf12), .B(_2264__bF_buf2), .C(regs_0__20_), .Y(_2386_) );
OAI21X1 OAI21X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf4), .B(_1041__bF_buf0), .C(_2386_), .Y(_12_) );
OAI21X1 OAI21X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf11), .B(_2264__bF_buf1), .C(regs_0__21_), .Y(_2387_) );
OAI21X1 OAI21X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf3), .B(_1043__bF_buf0), .C(_2387_), .Y(_13_) );
OAI21X1 OAI21X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf10), .B(_2264__bF_buf0), .C(regs_0__22_), .Y(_2388_) );
OAI21X1 OAI21X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf2), .B(_1045__bF_buf0), .C(_2388_), .Y(_14_) );
OAI21X1 OAI21X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf9), .B(_2264__bF_buf10), .C(regs_0__23_), .Y(_2389_) );
OAI21X1 OAI21X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf1), .B(_1047__bF_buf0), .C(_2389_), .Y(_15_) );
OAI21X1 OAI21X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf8), .B(_2264__bF_buf9), .C(regs_0__24_), .Y(_2390_) );
OAI21X1 OAI21X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf0), .B(_1049__bF_buf0), .C(_2390_), .Y(_16_) );
OAI21X1 OAI21X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf7), .B(_2264__bF_buf8), .C(regs_0__25_), .Y(_2391_) );
OAI21X1 OAI21X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf4), .B(_1051__bF_buf0), .C(_2391_), .Y(_17_) );
OAI21X1 OAI21X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf6), .B(_2264__bF_buf7), .C(regs_0__26_), .Y(_2392_) );
OAI21X1 OAI21X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf3), .B(_1053__bF_buf0), .C(_2392_), .Y(_18_) );
OAI21X1 OAI21X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf5), .B(_2264__bF_buf6), .C(regs_0__27_), .Y(_2393_) );
OAI21X1 OAI21X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf2), .B(_1055__bF_buf0), .C(_2393_), .Y(_19_) );
OAI21X1 OAI21X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf4), .B(_2264__bF_buf5), .C(regs_0__28_), .Y(_2394_) );
OAI21X1 OAI21X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf1), .B(_1057__bF_buf0), .C(_2394_), .Y(_20_) );
OAI21X1 OAI21X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf3), .B(_2264__bF_buf4), .C(regs_0__29_), .Y(_2395_) );
OAI21X1 OAI21X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf0), .B(_1059__bF_buf0), .C(_2395_), .Y(_21_) );
OAI21X1 OAI21X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf2), .B(_2264__bF_buf3), .C(regs_0__30_), .Y(_2396_) );
OAI21X1 OAI21X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf4), .B(_1061__bF_buf0), .C(_2396_), .Y(_23_) );
OAI21X1 OAI21X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf1), .B(_2264__bF_buf2), .C(regs_0__31_), .Y(_2397_) );
OAI21X1 OAI21X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_2365__bF_buf3), .B(_1063__bF_buf0), .C(_2397_), .Y(_24_) );
INVX8 INVX8_2 ( .gnd(gnd), .vdd(vdd), .A(raddr1[3]), .Y(_2398_) );
INVX8 INVX8_3 ( .gnd(gnd), .vdd(vdd), .A(raddr1_2_bF_buf10_), .Y(_2399_) );
NAND2X1 NAND2X1_298 ( .gnd(gnd), .vdd(vdd), .A(regs_22__0_), .B(raddr1_0_bF_buf96_), .Y(_2400_) );
OAI21X1 OAI21X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_1307_), .B(raddr1_0_bF_buf95_), .C(_2400_), .Y(_2401_) );
NAND2X1 NAND2X1_299 ( .gnd(gnd), .vdd(vdd), .A(regs_20__0_), .B(raddr1_0_bF_buf94_), .Y(_2402_) );
OAI21X1 OAI21X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_1407_), .B(raddr1_0_bF_buf93_), .C(_2402_), .Y(_2403_) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_2403_), .B(_2401_), .S(raddr1_1_bF_buf14_bF_buf3_), .Y(_2404_) );
NAND2X1 NAND2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf8), .B(_2404_), .Y(_2405_) );
NAND2X1 NAND2X1_301 ( .gnd(gnd), .vdd(vdd), .A(regs_18__0_), .B(raddr1_0_bF_buf92_), .Y(_2406_) );
OAI21X1 OAI21X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_1505_), .B(raddr1_0_bF_buf91_), .C(_2406_), .Y(_2407_) );
NAND2X1 NAND2X1_302 ( .gnd(gnd), .vdd(vdd), .A(regs_16__0_), .B(raddr1_0_bF_buf90_), .Y(_2408_) );
OAI21X1 OAI21X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_1604_), .B(raddr1_0_bF_buf89_), .C(_2408_), .Y(_2409_) );
MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_2409_), .B(_2407_), .S(raddr1_1_bF_buf13_bF_buf3_), .Y(_2410_) );
AOI21X1 AOI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(raddr1_2_bF_buf9_), .B(_2410_), .C(_2398__bF_buf7), .Y(_2411_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(regs_26__0_), .B(raddr1_0_bF_buf88_), .Y(_2412_) );
OAI21X1 OAI21X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_1138_), .B(raddr1_0_bF_buf87_), .C(raddr1_2_bF_buf8_), .Y(_2413_) );
NOR2X1 NOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_2412_), .B(_2413_), .Y(_2414_) );
INVX8 INVX8_4 ( .gnd(gnd), .vdd(vdd), .A(raddr1_1_bF_buf12_bF_buf3_), .Y(_2415_) );
OAI21X1 OAI21X1_1054 ( .gnd(gnd), .vdd(vdd), .A(regs_30__0_), .B(raddr1_2_bF_buf7_), .C(_2415__bF_buf8), .Y(_2416_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(regs_25__0_), .Y(_2417_) );
OAI21X1 OAI21X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_2417_), .B(raddr1_0_bF_buf86_), .C(raddr1_2_bF_buf6_), .Y(_2418_) );
AOI21X1 AOI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(regs_24__0_), .B(raddr1_0_bF_buf85_), .C(_2418_), .Y(_2419_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(regs_29__0_), .Y(_2420_) );
NOR2X1 NOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf84_), .B(_2420_), .Y(_2421_) );
NAND2X1 NAND2X1_303 ( .gnd(gnd), .vdd(vdd), .A(regs_28__0_), .B(raddr1_0_bF_buf83_), .Y(_2422_) );
NAND2X1 NAND2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf7), .B(_2422_), .Y(_2423_) );
OAI21X1 OAI21X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_2423_), .B(_2421_), .C(raddr1_1_bF_buf11_bF_buf3_), .Y(_2424_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_2414_), .B(_2416_), .C(_2424_), .D(_2419_), .Y(_2425_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_2425_), .B(_2398__bF_buf6), .C(_2405_), .D(_2411_), .Y(_2426_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(regs_5__0_), .Y(_2427_) );
OAI21X1 OAI21X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_2427_), .B(raddr1_0_bF_buf82_), .C(raddr1_1_bF_buf10_bF_buf3_), .Y(_2428_) );
AOI21X1 AOI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(regs_4__0_), .B(raddr1_0_bF_buf81_), .C(_2428_), .Y(_2429_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(regs_6__0_), .B(raddr1_0_bF_buf80_), .Y(_2430_) );
OAI21X1 OAI21X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_2097_), .B(raddr1_0_bF_buf79_), .C(_2415__bF_buf7), .Y(_2431_) );
OAI21X1 OAI21X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_2431_), .B(_2430_), .C(_2399__bF_buf6), .Y(_2432_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(regs_1__0_), .Y(_2433_) );
OAI21X1 OAI21X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_2433_), .B(raddr1_0_bF_buf78_), .C(raddr1_1_bF_buf9_bF_buf3_), .Y(_2434_) );
AOI21X1 AOI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(regs_0__0_), .B(raddr1_0_bF_buf77_), .C(_2434_), .Y(_2435_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(regs_3__0_), .Y(_2436_) );
AOI21X1 AOI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(regs_2__0_), .B(raddr1_0_bF_buf76_), .C(raddr1_1_bF_buf8_), .Y(_2437_) );
OAI21X1 OAI21X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_2436_), .B(raddr1_0_bF_buf75_), .C(_2437_), .Y(_2438_) );
NAND2X1 NAND2X1_305 ( .gnd(gnd), .vdd(vdd), .A(raddr1_2_bF_buf5_), .B(_2438_), .Y(_2439_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_2439_), .B(_2435_), .C(_2432_), .D(_2429_), .Y(_2440_) );
NAND2X1 NAND2X1_306 ( .gnd(gnd), .vdd(vdd), .A(regs_10__0_), .B(raddr1_0_bF_buf74_), .Y(_2441_) );
OAI21X1 OAI21X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_1900_), .B(raddr1_0_bF_buf73_), .C(_2441_), .Y(_2442_) );
NAND2X1 NAND2X1_307 ( .gnd(gnd), .vdd(vdd), .A(regs_8__0_), .B(raddr1_0_bF_buf72_), .Y(_2443_) );
OAI21X1 OAI21X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_1999_), .B(raddr1_0_bF_buf71_), .C(_2443_), .Y(_2444_) );
MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_2444_), .B(_2442_), .S(raddr1_1_bF_buf7_), .Y(_2445_) );
NAND2X1 NAND2X1_308 ( .gnd(gnd), .vdd(vdd), .A(regs_14__0_), .B(raddr1_0_bF_buf70_), .Y(_2446_) );
OAI21X1 OAI21X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_1702_), .B(raddr1_0_bF_buf69_), .C(_2446_), .Y(_2447_) );
NAND2X1 NAND2X1_309 ( .gnd(gnd), .vdd(vdd), .A(regs_12__0_), .B(raddr1_0_bF_buf68_), .Y(_2448_) );
OAI21X1 OAI21X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_1802_), .B(raddr1_0_bF_buf67_), .C(_2448_), .Y(_2449_) );
MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_2449_), .B(_2447_), .S(raddr1_1_bF_buf6_), .Y(_2450_) );
MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_2450_), .B(_2445_), .S(_2399__bF_buf5), .Y(_2451_) );
MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_2451_), .B(_2440_), .S(_2398__bF_buf5), .Y(_2452_) );
MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_2452_), .B(_2426_), .S(raddr1_4_bF_buf4_), .Y(_5511__0_) );
OAI21X1 OAI21X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_1410_), .B(raddr1_0_bF_buf66_), .C(raddr1_1_bF_buf5_), .Y(_2453_) );
AOI21X1 AOI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(regs_20__1_), .B(raddr1_0_bF_buf65_), .C(_2453_), .Y(_2454_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(regs_22__1_), .B(raddr1_0_bF_buf64_), .Y(_2455_) );
OAI21X1 OAI21X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_1312_), .B(raddr1_0_bF_buf63_), .C(_2415__bF_buf6), .Y(_2456_) );
OAI21X1 OAI21X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_2456_), .B(_2455_), .C(_2399__bF_buf4), .Y(_2457_) );
OAI21X1 OAI21X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_1607_), .B(raddr1_0_bF_buf62_), .C(raddr1_1_bF_buf4_), .Y(_2458_) );
AOI21X1 AOI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(regs_16__1_), .B(raddr1_0_bF_buf61_), .C(_2458_), .Y(_2459_) );
NOR2X1 NOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf60_), .B(_1509_), .Y(_2460_) );
NAND2X1 NAND2X1_310 ( .gnd(gnd), .vdd(vdd), .A(regs_18__1_), .B(raddr1_0_bF_buf59_), .Y(_2461_) );
NAND2X1 NAND2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf5), .B(_2461_), .Y(_2462_) );
OAI21X1 OAI21X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_2462_), .B(_2460_), .C(raddr1_2_bF_buf4_), .Y(_2463_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_2459_), .B(_2463_), .C(_2457_), .D(_2454_), .Y(_2464_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(regs_29__1_), .Y(_2465_) );
NAND2X1 NAND2X1_312 ( .gnd(gnd), .vdd(vdd), .A(regs_28__1_), .B(raddr1_0_bF_buf58_), .Y(_2466_) );
OAI21X1 OAI21X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_2465_), .B(raddr1_0_bF_buf57_), .C(_2466_), .Y(_2467_) );
MUX2X1 MUX2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_2467_), .B(regs_30__1_), .S(raddr1_1_bF_buf3_), .Y(_2468_) );
NAND2X1 NAND2X1_313 ( .gnd(gnd), .vdd(vdd), .A(regs_26__1_), .B(raddr1_0_bF_buf56_), .Y(_2469_) );
OAI21X1 OAI21X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_1145_), .B(raddr1_0_bF_buf55_), .C(_2469_), .Y(_2470_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(regs_25__1_), .Y(_2471_) );
NAND2X1 NAND2X1_314 ( .gnd(gnd), .vdd(vdd), .A(regs_24__1_), .B(raddr1_0_bF_buf54_), .Y(_2472_) );
OAI21X1 OAI21X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_2471_), .B(raddr1_0_bF_buf53_), .C(_2472_), .Y(_2473_) );
MUX2X1 MUX2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_2473_), .B(_2470_), .S(raddr1_1_bF_buf2_), .Y(_2474_) );
MUX2X1 MUX2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_2474_), .B(_2468_), .S(raddr1_2_bF_buf3_), .Y(_2475_) );
MUX2X1 MUX2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_2475_), .B(_2464_), .S(_2398__bF_buf4), .Y(_2476_) );
NAND2X1 NAND2X1_315 ( .gnd(gnd), .vdd(vdd), .A(regs_6__1_), .B(raddr1_0_bF_buf52_), .Y(_2477_) );
OAI21X1 OAI21X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_2103_), .B(raddr1_0_bF_buf51_), .C(_2477_), .Y(_2478_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(regs_5__1_), .Y(_2479_) );
NAND2X1 NAND2X1_316 ( .gnd(gnd), .vdd(vdd), .A(regs_4__1_), .B(raddr1_0_bF_buf50_), .Y(_2480_) );
OAI21X1 OAI21X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_2479_), .B(raddr1_0_bF_buf49_), .C(_2480_), .Y(_2481_) );
MUX2X1 MUX2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_2481_), .B(_2478_), .S(raddr1_1_bF_buf1_), .Y(_2482_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(regs_3__1_), .Y(_2483_) );
NAND2X1 NAND2X1_317 ( .gnd(gnd), .vdd(vdd), .A(regs_2__1_), .B(raddr1_0_bF_buf48_), .Y(_2484_) );
OAI21X1 OAI21X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_2483_), .B(raddr1_0_bF_buf47_), .C(_2484_), .Y(_2485_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(regs_1__1_), .Y(_2486_) );
NAND2X1 NAND2X1_318 ( .gnd(gnd), .vdd(vdd), .A(regs_0__1_), .B(raddr1_0_bF_buf46_), .Y(_2487_) );
OAI21X1 OAI21X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_2486_), .B(raddr1_0_bF_buf45_), .C(_2487_), .Y(_2488_) );
MUX2X1 MUX2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_2488_), .B(_2485_), .S(raddr1_1_bF_buf0_), .Y(_2489_) );
MUX2X1 MUX2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_2489_), .B(_2482_), .S(raddr1_2_bF_buf2_), .Y(_2490_) );
NAND2X1 NAND2X1_319 ( .gnd(gnd), .vdd(vdd), .A(regs_10__1_), .B(raddr1_0_bF_buf44_), .Y(_2491_) );
OAI21X1 OAI21X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_1904_), .B(raddr1_0_bF_buf43_), .C(_2491_), .Y(_2492_) );
NAND2X1 NAND2X1_320 ( .gnd(gnd), .vdd(vdd), .A(regs_8__1_), .B(raddr1_0_bF_buf42_), .Y(_2493_) );
OAI21X1 OAI21X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_2002_), .B(raddr1_0_bF_buf41_), .C(_2493_), .Y(_2494_) );
MUX2X1 MUX2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_2494_), .B(_2492_), .S(raddr1_1_bF_buf14_bF_buf2_), .Y(_2495_) );
NAND2X1 NAND2X1_321 ( .gnd(gnd), .vdd(vdd), .A(regs_14__1_), .B(raddr1_0_bF_buf40_), .Y(_2496_) );
OAI21X1 OAI21X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_1707_), .B(raddr1_0_bF_buf39_), .C(_2496_), .Y(_2497_) );
NAND2X1 NAND2X1_322 ( .gnd(gnd), .vdd(vdd), .A(regs_12__1_), .B(raddr1_0_bF_buf38_), .Y(_2498_) );
OAI21X1 OAI21X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_1805_), .B(raddr1_0_bF_buf37_), .C(_2498_), .Y(_2499_) );
MUX2X1 MUX2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_2499_), .B(_2497_), .S(raddr1_1_bF_buf13_bF_buf2_), .Y(_2500_) );
MUX2X1 MUX2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_2500_), .B(_2495_), .S(_2399__bF_buf3), .Y(_2501_) );
MUX2X1 MUX2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_2501_), .B(_2490_), .S(_2398__bF_buf3), .Y(_2502_) );
MUX2X1 MUX2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_2502_), .B(_2476_), .S(raddr1_4_bF_buf3_), .Y(_5511__1_) );
NAND2X1 NAND2X1_323 ( .gnd(gnd), .vdd(vdd), .A(regs_22__2_), .B(raddr1_0_bF_buf36_), .Y(_2503_) );
OAI21X1 OAI21X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_1314_), .B(raddr1_0_bF_buf35_), .C(_2503_), .Y(_2504_) );
NAND2X1 NAND2X1_324 ( .gnd(gnd), .vdd(vdd), .A(regs_20__2_), .B(raddr1_0_bF_buf34_), .Y(_2505_) );
OAI21X1 OAI21X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_1412_), .B(raddr1_0_bF_buf33_), .C(_2505_), .Y(_2506_) );
MUX2X1 MUX2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_2506_), .B(_2504_), .S(raddr1_1_bF_buf12_bF_buf2_), .Y(_2507_) );
NAND2X1 NAND2X1_325 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf2), .B(_2507_), .Y(_2508_) );
NAND2X1 NAND2X1_326 ( .gnd(gnd), .vdd(vdd), .A(regs_18__2_), .B(raddr1_0_bF_buf32_), .Y(_2509_) );
OAI21X1 OAI21X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_1511_), .B(raddr1_0_bF_buf31_), .C(_2509_), .Y(_2510_) );
NAND2X1 NAND2X1_327 ( .gnd(gnd), .vdd(vdd), .A(regs_16__2_), .B(raddr1_0_bF_buf30_), .Y(_2511_) );
OAI21X1 OAI21X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_1609_), .B(raddr1_0_bF_buf29_), .C(_2511_), .Y(_2512_) );
MUX2X1 MUX2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_2512_), .B(_2510_), .S(raddr1_1_bF_buf11_bF_buf2_), .Y(_2513_) );
AOI21X1 AOI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(raddr1_2_bF_buf1_), .B(_2513_), .C(_2398__bF_buf2), .Y(_2514_) );
OAI21X1 OAI21X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_1147_), .B(raddr1_0_bF_buf28_), .C(raddr1_2_bF_buf0_), .Y(_2515_) );
AOI21X1 AOI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(regs_26__2_), .B(raddr1_0_bF_buf27_), .C(_2515_), .Y(_2516_) );
OAI21X1 OAI21X1_1087 ( .gnd(gnd), .vdd(vdd), .A(regs_30__2_), .B(raddr1_2_bF_buf10_), .C(_2415__bF_buf4), .Y(_2517_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(regs_25__2_), .Y(_2518_) );
OAI21X1 OAI21X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_2518_), .B(raddr1_0_bF_buf26_), .C(raddr1_2_bF_buf9_), .Y(_2519_) );
AOI21X1 AOI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(regs_24__2_), .B(raddr1_0_bF_buf25_), .C(_2519_), .Y(_2520_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(regs_29__2_), .Y(_2521_) );
NOR2X1 NOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf24_), .B(_2521_), .Y(_2522_) );
NAND2X1 NAND2X1_328 ( .gnd(gnd), .vdd(vdd), .A(regs_28__2_), .B(raddr1_0_bF_buf23_), .Y(_2523_) );
NAND2X1 NAND2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf1), .B(_2523_), .Y(_2524_) );
OAI21X1 OAI21X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_2524_), .B(_2522_), .C(raddr1_1_bF_buf10_bF_buf2_), .Y(_2525_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_2516_), .B(_2517_), .C(_2525_), .D(_2520_), .Y(_2526_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_2526_), .B(_2398__bF_buf1), .C(_2508_), .D(_2514_), .Y(_2527_) );
NAND2X1 NAND2X1_330 ( .gnd(gnd), .vdd(vdd), .A(regs_6__2_), .B(raddr1_0_bF_buf22_), .Y(_2528_) );
OAI21X1 OAI21X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_2105_), .B(raddr1_0_bF_buf21_), .C(_2528_), .Y(_2529_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(regs_5__2_), .Y(_2530_) );
NAND2X1 NAND2X1_331 ( .gnd(gnd), .vdd(vdd), .A(regs_4__2_), .B(raddr1_0_bF_buf20_), .Y(_2531_) );
OAI21X1 OAI21X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_2530_), .B(raddr1_0_bF_buf19_), .C(_2531_), .Y(_2532_) );
MUX2X1 MUX2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_2532_), .B(_2529_), .S(raddr1_1_bF_buf9_bF_buf2_), .Y(_2533_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(regs_3__2_), .Y(_2534_) );
NAND2X1 NAND2X1_332 ( .gnd(gnd), .vdd(vdd), .A(regs_2__2_), .B(raddr1_0_bF_buf18_), .Y(_2535_) );
OAI21X1 OAI21X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_2534_), .B(raddr1_0_bF_buf17_), .C(_2535_), .Y(_2536_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(regs_1__2_), .Y(_2537_) );
NAND2X1 NAND2X1_333 ( .gnd(gnd), .vdd(vdd), .A(regs_0__2_), .B(raddr1_0_bF_buf16_), .Y(_2538_) );
OAI21X1 OAI21X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_2537_), .B(raddr1_0_bF_buf15_), .C(_2538_), .Y(_2539_) );
MUX2X1 MUX2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_2539_), .B(_2536_), .S(raddr1_1_bF_buf8_), .Y(_2540_) );
MUX2X1 MUX2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_2540_), .B(_2533_), .S(raddr1_2_bF_buf8_), .Y(_2541_) );
NAND2X1 NAND2X1_334 ( .gnd(gnd), .vdd(vdd), .A(regs_14__2_), .B(raddr1_0_bF_buf14_), .Y(_2542_) );
OAI21X1 OAI21X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_1709_), .B(raddr1_0_bF_buf13_), .C(_2542_), .Y(_2543_) );
NAND2X1 NAND2X1_335 ( .gnd(gnd), .vdd(vdd), .A(regs_12__2_), .B(raddr1_0_bF_buf12_), .Y(_2544_) );
OAI21X1 OAI21X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_1807_), .B(raddr1_0_bF_buf11_), .C(_2544_), .Y(_2545_) );
MUX2X1 MUX2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_2545_), .B(_2543_), .S(raddr1_1_bF_buf7_), .Y(_2546_) );
NAND2X1 NAND2X1_336 ( .gnd(gnd), .vdd(vdd), .A(regs_10__2_), .B(raddr1_0_bF_buf10_), .Y(_2547_) );
OAI21X1 OAI21X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_1906_), .B(raddr1_0_bF_buf9_), .C(_2547_), .Y(_2548_) );
NAND2X1 NAND2X1_337 ( .gnd(gnd), .vdd(vdd), .A(regs_8__2_), .B(raddr1_0_bF_buf8_), .Y(_2549_) );
OAI21X1 OAI21X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_2004_), .B(raddr1_0_bF_buf7_), .C(_2549_), .Y(_2550_) );
MUX2X1 MUX2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_2550_), .B(_2548_), .S(raddr1_1_bF_buf6_), .Y(_2551_) );
MUX2X1 MUX2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_2546_), .S(raddr1_2_bF_buf7_), .Y(_2552_) );
MUX2X1 MUX2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_2552_), .B(_2541_), .S(_2398__bF_buf0), .Y(_2553_) );
MUX2X1 MUX2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_2553_), .B(_2527_), .S(raddr1_4_bF_buf2_), .Y(_5511__2_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(regs_5__3_), .Y(_2554_) );
OAI21X1 OAI21X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_2554_), .B(raddr1_0_bF_buf6_), .C(raddr1_1_bF_buf5_), .Y(_2555_) );
AOI21X1 AOI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(regs_4__3_), .B(raddr1_0_bF_buf5_), .C(_2555_), .Y(_2556_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(regs_6__3_), .B(raddr1_0_bF_buf4_), .Y(_2557_) );
OAI21X1 OAI21X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_2107_), .B(raddr1_0_bF_buf3_), .C(_2415__bF_buf3), .Y(_2558_) );
OAI21X1 OAI21X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_2558_), .B(_2557_), .C(_2399__bF_buf0), .Y(_2559_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(regs_1__3_), .Y(_2560_) );
OAI21X1 OAI21X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_2560_), .B(raddr1_0_bF_buf2_), .C(raddr1_1_bF_buf4_), .Y(_2561_) );
AOI21X1 AOI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(regs_0__3_), .B(raddr1_0_bF_buf1_), .C(_2561_), .Y(_2562_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(regs_3__3_), .Y(_2563_) );
NOR2X1 NOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf0_), .B(_2563_), .Y(_2564_) );
NAND2X1 NAND2X1_338 ( .gnd(gnd), .vdd(vdd), .A(regs_2__3_), .B(raddr1_0_bF_buf96_), .Y(_2565_) );
NAND2X1 NAND2X1_339 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf2), .B(_2565_), .Y(_2566_) );
OAI21X1 OAI21X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_2566_), .B(_2564_), .C(raddr1_2_bF_buf6_), .Y(_2567_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_2562_), .B(_2567_), .C(_2559_), .D(_2556_), .Y(_2568_) );
NAND2X1 NAND2X1_340 ( .gnd(gnd), .vdd(vdd), .A(regs_10__3_), .B(raddr1_0_bF_buf95_), .Y(_2569_) );
OAI21X1 OAI21X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_1908_), .B(raddr1_0_bF_buf94_), .C(_2569_), .Y(_2570_) );
NAND2X1 NAND2X1_341 ( .gnd(gnd), .vdd(vdd), .A(regs_8__3_), .B(raddr1_0_bF_buf93_), .Y(_2571_) );
OAI21X1 OAI21X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .B(raddr1_0_bF_buf92_), .C(_2571_), .Y(_2572_) );
MUX2X1 MUX2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_2572_), .B(_2570_), .S(raddr1_1_bF_buf3_), .Y(_2573_) );
NAND2X1 NAND2X1_342 ( .gnd(gnd), .vdd(vdd), .A(regs_14__3_), .B(raddr1_0_bF_buf91_), .Y(_2574_) );
OAI21X1 OAI21X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_1711_), .B(raddr1_0_bF_buf90_), .C(_2574_), .Y(_2575_) );
NAND2X1 NAND2X1_343 ( .gnd(gnd), .vdd(vdd), .A(regs_12__3_), .B(raddr1_0_bF_buf89_), .Y(_2576_) );
OAI21X1 OAI21X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_1809_), .B(raddr1_0_bF_buf88_), .C(_2576_), .Y(_2577_) );
MUX2X1 MUX2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_2577_), .B(_2575_), .S(raddr1_1_bF_buf2_), .Y(_2578_) );
MUX2X1 MUX2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_2578_), .B(_2573_), .S(_2399__bF_buf8), .Y(_2579_) );
MUX2X1 MUX2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_2579_), .B(_2568_), .S(_2398__bF_buf7), .Y(_2580_) );
OAI21X1 OAI21X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_1611_), .B(raddr1_0_bF_buf87_), .C(raddr1_1_bF_buf1_), .Y(_2581_) );
AOI21X1 AOI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(regs_16__3_), .B(raddr1_0_bF_buf86_), .C(_2581_), .Y(_2582_) );
NOR2X1 NOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf85_), .B(_1513_), .Y(_2583_) );
NAND2X1 NAND2X1_344 ( .gnd(gnd), .vdd(vdd), .A(regs_18__3_), .B(raddr1_0_bF_buf84_), .Y(_2584_) );
NAND2X1 NAND2X1_345 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf1), .B(_2584_), .Y(_2585_) );
OAI21X1 OAI21X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_2585_), .B(_2583_), .C(raddr1_2_bF_buf5_), .Y(_2586_) );
OAI21X1 OAI21X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_1414_), .B(raddr1_0_bF_buf83_), .C(raddr1_1_bF_buf0_), .Y(_2587_) );
AOI21X1 AOI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(regs_20__3_), .B(raddr1_0_bF_buf82_), .C(_2587_), .Y(_2588_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(regs_22__3_), .B(raddr1_0_bF_buf81_), .Y(_2589_) );
OAI21X1 OAI21X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_1316_), .B(raddr1_0_bF_buf80_), .C(_2415__bF_buf0), .Y(_2590_) );
OAI21X1 OAI21X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .B(_2589_), .C(_2399__bF_buf7), .Y(_2591_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_2582_), .B(_2586_), .C(_2591_), .D(_2588_), .Y(_2592_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(regs_29__3_), .Y(_2593_) );
NAND2X1 NAND2X1_346 ( .gnd(gnd), .vdd(vdd), .A(regs_28__3_), .B(raddr1_0_bF_buf79_), .Y(_2594_) );
OAI21X1 OAI21X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_2593_), .B(raddr1_0_bF_buf78_), .C(_2594_), .Y(_2595_) );
MUX2X1 MUX2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_2595_), .B(regs_30__3_), .S(raddr1_1_bF_buf14_bF_buf1_), .Y(_2596_) );
NAND2X1 NAND2X1_347 ( .gnd(gnd), .vdd(vdd), .A(regs_26__3_), .B(raddr1_0_bF_buf77_), .Y(_2597_) );
OAI21X1 OAI21X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_1149_), .B(raddr1_0_bF_buf76_), .C(_2597_), .Y(_2598_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(regs_25__3_), .Y(_2599_) );
NAND2X1 NAND2X1_348 ( .gnd(gnd), .vdd(vdd), .A(regs_24__3_), .B(raddr1_0_bF_buf75_), .Y(_2600_) );
OAI21X1 OAI21X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_2599_), .B(raddr1_0_bF_buf74_), .C(_2600_), .Y(_2601_) );
MUX2X1 MUX2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_2601_), .B(_2598_), .S(raddr1_1_bF_buf13_bF_buf1_), .Y(_2602_) );
MUX2X1 MUX2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_2602_), .B(_2596_), .S(raddr1_2_bF_buf4_), .Y(_2603_) );
MUX2X1 MUX2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_2603_), .B(_2592_), .S(_2398__bF_buf6), .Y(_2604_) );
MUX2X1 MUX2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_2580_), .B(_2604_), .S(raddr1_4_bF_buf1_), .Y(_5511__3_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(regs_5__4_), .Y(_2605_) );
OAI21X1 OAI21X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_2605_), .B(raddr1_0_bF_buf73_), .C(raddr1_1_bF_buf12_bF_buf1_), .Y(_2606_) );
AOI21X1 AOI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(regs_4__4_), .B(raddr1_0_bF_buf72_), .C(_2606_), .Y(_2607_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(regs_6__4_), .B(raddr1_0_bF_buf71_), .Y(_2608_) );
OAI21X1 OAI21X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_2109_), .B(raddr1_0_bF_buf70_), .C(_2415__bF_buf8), .Y(_2609_) );
OAI21X1 OAI21X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_2609_), .B(_2608_), .C(_2399__bF_buf6), .Y(_2610_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(regs_1__4_), .Y(_2611_) );
OAI21X1 OAI21X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_2611_), .B(raddr1_0_bF_buf69_), .C(raddr1_1_bF_buf11_bF_buf1_), .Y(_2612_) );
AOI21X1 AOI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(regs_0__4_), .B(raddr1_0_bF_buf68_), .C(_2612_), .Y(_2613_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(regs_3__4_), .Y(_2614_) );
NOR2X1 NOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf67_), .B(_2614_), .Y(_2615_) );
NAND2X1 NAND2X1_349 ( .gnd(gnd), .vdd(vdd), .A(regs_2__4_), .B(raddr1_0_bF_buf66_), .Y(_2616_) );
NAND2X1 NAND2X1_350 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf7), .B(_2616_), .Y(_2617_) );
OAI21X1 OAI21X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_2617_), .B(_2615_), .C(raddr1_2_bF_buf3_), .Y(_2618_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_2613_), .B(_2618_), .C(_2610_), .D(_2607_), .Y(_2619_) );
NAND2X1 NAND2X1_351 ( .gnd(gnd), .vdd(vdd), .A(regs_10__4_), .B(raddr1_0_bF_buf65_), .Y(_2620_) );
OAI21X1 OAI21X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_1910_), .B(raddr1_0_bF_buf64_), .C(_2620_), .Y(_2621_) );
NAND2X1 NAND2X1_352 ( .gnd(gnd), .vdd(vdd), .A(regs_8__4_), .B(raddr1_0_bF_buf63_), .Y(_2622_) );
OAI21X1 OAI21X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_2008_), .B(raddr1_0_bF_buf62_), .C(_2622_), .Y(_2623_) );
MUX2X1 MUX2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_2623_), .B(_2621_), .S(raddr1_1_bF_buf10_bF_buf1_), .Y(_2624_) );
NAND2X1 NAND2X1_353 ( .gnd(gnd), .vdd(vdd), .A(regs_14__4_), .B(raddr1_0_bF_buf61_), .Y(_2625_) );
OAI21X1 OAI21X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_1713_), .B(raddr1_0_bF_buf60_), .C(_2625_), .Y(_2626_) );
NAND2X1 NAND2X1_354 ( .gnd(gnd), .vdd(vdd), .A(regs_12__4_), .B(raddr1_0_bF_buf59_), .Y(_2627_) );
OAI21X1 OAI21X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_1811_), .B(raddr1_0_bF_buf58_), .C(_2627_), .Y(_2628_) );
MUX2X1 MUX2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_2628_), .B(_2626_), .S(raddr1_1_bF_buf9_bF_buf1_), .Y(_2629_) );
MUX2X1 MUX2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_2629_), .B(_2624_), .S(_2399__bF_buf5), .Y(_2630_) );
MUX2X1 MUX2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_2630_), .B(_2619_), .S(_2398__bF_buf5), .Y(_2631_) );
OAI21X1 OAI21X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_1613_), .B(raddr1_0_bF_buf57_), .C(raddr1_1_bF_buf8_), .Y(_2632_) );
AOI21X1 AOI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(regs_16__4_), .B(raddr1_0_bF_buf56_), .C(_2632_), .Y(_2633_) );
NOR2X1 NOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf55_), .B(_1515_), .Y(_2634_) );
NAND2X1 NAND2X1_355 ( .gnd(gnd), .vdd(vdd), .A(regs_18__4_), .B(raddr1_0_bF_buf54_), .Y(_2635_) );
NAND2X1 NAND2X1_356 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf6), .B(_2635_), .Y(_2636_) );
OAI21X1 OAI21X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_2636_), .B(_2634_), .C(raddr1_2_bF_buf2_), .Y(_2637_) );
OAI21X1 OAI21X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_1416_), .B(raddr1_0_bF_buf53_), .C(raddr1_1_bF_buf7_), .Y(_2638_) );
AOI21X1 AOI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(regs_20__4_), .B(raddr1_0_bF_buf52_), .C(_2638_), .Y(_2639_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(regs_22__4_), .B(raddr1_0_bF_buf51_), .Y(_2640_) );
OAI21X1 OAI21X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_1318_), .B(raddr1_0_bF_buf50_), .C(_2415__bF_buf5), .Y(_2641_) );
OAI21X1 OAI21X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_2641_), .B(_2640_), .C(_2399__bF_buf4), .Y(_2642_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_2633_), .B(_2637_), .C(_2642_), .D(_2639_), .Y(_2643_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(regs_29__4_), .Y(_2644_) );
NAND2X1 NAND2X1_357 ( .gnd(gnd), .vdd(vdd), .A(regs_28__4_), .B(raddr1_0_bF_buf49_), .Y(_2645_) );
OAI21X1 OAI21X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_2644_), .B(raddr1_0_bF_buf48_), .C(_2645_), .Y(_2646_) );
MUX2X1 MUX2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_2646_), .B(regs_30__4_), .S(raddr1_1_bF_buf6_), .Y(_2647_) );
NAND2X1 NAND2X1_358 ( .gnd(gnd), .vdd(vdd), .A(regs_26__4_), .B(raddr1_0_bF_buf47_), .Y(_2648_) );
OAI21X1 OAI21X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_1151_), .B(raddr1_0_bF_buf46_), .C(_2648_), .Y(_2649_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(regs_25__4_), .Y(_2650_) );
NAND2X1 NAND2X1_359 ( .gnd(gnd), .vdd(vdd), .A(regs_24__4_), .B(raddr1_0_bF_buf45_), .Y(_2651_) );
OAI21X1 OAI21X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_2650_), .B(raddr1_0_bF_buf44_), .C(_2651_), .Y(_2652_) );
MUX2X1 MUX2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_2652_), .B(_2649_), .S(raddr1_1_bF_buf5_), .Y(_2653_) );
MUX2X1 MUX2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_2653_), .B(_2647_), .S(raddr1_2_bF_buf1_), .Y(_2654_) );
MUX2X1 MUX2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_2654_), .B(_2643_), .S(_2398__bF_buf4), .Y(_2655_) );
MUX2X1 MUX2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_2631_), .B(_2655_), .S(raddr1_4_bF_buf0_), .Y(_5511__4_) );
OAI21X1 OAI21X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_1418_), .B(raddr1_0_bF_buf43_), .C(raddr1_1_bF_buf4_), .Y(_2656_) );
AOI21X1 AOI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(regs_20__5_), .B(raddr1_0_bF_buf42_), .C(_2656_), .Y(_2657_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(regs_22__5_), .B(raddr1_0_bF_buf41_), .Y(_2658_) );
OAI21X1 OAI21X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_1320_), .B(raddr1_0_bF_buf40_), .C(_2415__bF_buf4), .Y(_2659_) );
OAI21X1 OAI21X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_2659_), .B(_2658_), .C(_2399__bF_buf3), .Y(_2660_) );
OAI21X1 OAI21X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(raddr1_0_bF_buf39_), .C(raddr1_1_bF_buf3_), .Y(_2661_) );
AOI21X1 AOI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(regs_16__5_), .B(raddr1_0_bF_buf38_), .C(_2661_), .Y(_2662_) );
NOR2X1 NOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf37_), .B(_1517_), .Y(_2663_) );
NAND2X1 NAND2X1_360 ( .gnd(gnd), .vdd(vdd), .A(regs_18__5_), .B(raddr1_0_bF_buf36_), .Y(_2664_) );
NAND2X1 NAND2X1_361 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf3), .B(_2664_), .Y(_2665_) );
OAI21X1 OAI21X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_2665_), .B(_2663_), .C(raddr1_2_bF_buf0_), .Y(_2666_) );
OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_2662_), .B(_2666_), .C(_2660_), .D(_2657_), .Y(_2667_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(regs_29__5_), .Y(_2668_) );
NAND2X1 NAND2X1_362 ( .gnd(gnd), .vdd(vdd), .A(regs_28__5_), .B(raddr1_0_bF_buf35_), .Y(_2669_) );
OAI21X1 OAI21X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_2668_), .B(raddr1_0_bF_buf34_), .C(_2669_), .Y(_2670_) );
MUX2X1 MUX2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_2670_), .B(regs_30__5_), .S(raddr1_1_bF_buf2_), .Y(_2671_) );
NAND2X1 NAND2X1_363 ( .gnd(gnd), .vdd(vdd), .A(regs_26__5_), .B(raddr1_0_bF_buf33_), .Y(_2672_) );
OAI21X1 OAI21X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(raddr1_0_bF_buf32_), .C(_2672_), .Y(_2673_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(regs_25__5_), .Y(_2674_) );
NAND2X1 NAND2X1_364 ( .gnd(gnd), .vdd(vdd), .A(regs_24__5_), .B(raddr1_0_bF_buf31_), .Y(_2675_) );
OAI21X1 OAI21X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_2674_), .B(raddr1_0_bF_buf30_), .C(_2675_), .Y(_2676_) );
MUX2X1 MUX2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_2676_), .B(_2673_), .S(raddr1_1_bF_buf1_), .Y(_2677_) );
MUX2X1 MUX2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_2677_), .B(_2671_), .S(raddr1_2_bF_buf10_), .Y(_2678_) );
MUX2X1 MUX2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_2678_), .B(_2667_), .S(_2398__bF_buf3), .Y(_2679_) );
NAND2X1 NAND2X1_365 ( .gnd(gnd), .vdd(vdd), .A(regs_6__5_), .B(raddr1_0_bF_buf29_), .Y(_2680_) );
OAI21X1 OAI21X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_2111_), .B(raddr1_0_bF_buf28_), .C(_2680_), .Y(_2681_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(regs_5__5_), .Y(_2682_) );
NAND2X1 NAND2X1_366 ( .gnd(gnd), .vdd(vdd), .A(regs_4__5_), .B(raddr1_0_bF_buf27_), .Y(_2683_) );
OAI21X1 OAI21X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_2682_), .B(raddr1_0_bF_buf26_), .C(_2683_), .Y(_2684_) );
MUX2X1 MUX2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_2684_), .B(_2681_), .S(raddr1_1_bF_buf0_), .Y(_2685_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(regs_3__5_), .Y(_2686_) );
NAND2X1 NAND2X1_367 ( .gnd(gnd), .vdd(vdd), .A(regs_2__5_), .B(raddr1_0_bF_buf25_), .Y(_2687_) );
OAI21X1 OAI21X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_2686_), .B(raddr1_0_bF_buf24_), .C(_2687_), .Y(_2688_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(regs_1__5_), .Y(_2689_) );
NAND2X1 NAND2X1_368 ( .gnd(gnd), .vdd(vdd), .A(regs_0__5_), .B(raddr1_0_bF_buf23_), .Y(_2690_) );
OAI21X1 OAI21X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_2689_), .B(raddr1_0_bF_buf22_), .C(_2690_), .Y(_2691_) );
MUX2X1 MUX2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_2691_), .B(_2688_), .S(raddr1_1_bF_buf14_bF_buf0_), .Y(_2692_) );
MUX2X1 MUX2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_2692_), .B(_2685_), .S(raddr1_2_bF_buf9_), .Y(_2693_) );
NAND2X1 NAND2X1_369 ( .gnd(gnd), .vdd(vdd), .A(regs_14__5_), .B(raddr1_0_bF_buf21_), .Y(_2694_) );
OAI21X1 OAI21X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_1715_), .B(raddr1_0_bF_buf20_), .C(_2694_), .Y(_2695_) );
NAND2X1 NAND2X1_370 ( .gnd(gnd), .vdd(vdd), .A(regs_12__5_), .B(raddr1_0_bF_buf19_), .Y(_2696_) );
OAI21X1 OAI21X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_1813_), .B(raddr1_0_bF_buf18_), .C(_2696_), .Y(_2697_) );
MUX2X1 MUX2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_2697_), .B(_2695_), .S(raddr1_1_bF_buf13_bF_buf0_), .Y(_2698_) );
NAND2X1 NAND2X1_371 ( .gnd(gnd), .vdd(vdd), .A(regs_10__5_), .B(raddr1_0_bF_buf17_), .Y(_2699_) );
OAI21X1 OAI21X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_1912_), .B(raddr1_0_bF_buf16_), .C(_2699_), .Y(_2700_) );
NAND2X1 NAND2X1_372 ( .gnd(gnd), .vdd(vdd), .A(regs_8__5_), .B(raddr1_0_bF_buf15_), .Y(_2701_) );
OAI21X1 OAI21X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_2010_), .B(raddr1_0_bF_buf14_), .C(_2701_), .Y(_2702_) );
MUX2X1 MUX2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_2702_), .B(_2700_), .S(raddr1_1_bF_buf12_bF_buf0_), .Y(_2703_) );
MUX2X1 MUX2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_2703_), .B(_2698_), .S(raddr1_2_bF_buf8_), .Y(_2704_) );
MUX2X1 MUX2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_2704_), .B(_2693_), .S(_2398__bF_buf2), .Y(_2705_) );
MUX2X1 MUX2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_2705_), .B(_2679_), .S(raddr1_4_bF_buf4_), .Y(_5511__5_) );
OAI21X1 OAI21X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(raddr1_0_bF_buf13_), .C(raddr1_1_bF_buf11_bF_buf0_), .Y(_2706_) );
AOI21X1 AOI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(regs_20__6_), .B(raddr1_0_bF_buf12_), .C(_2706_), .Y(_2707_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(regs_22__6_), .B(raddr1_0_bF_buf11_), .Y(_2708_) );
OAI21X1 OAI21X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_1322_), .B(raddr1_0_bF_buf10_), .C(_2415__bF_buf2), .Y(_2709_) );
OAI21X1 OAI21X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_2709_), .B(_2708_), .C(_2399__bF_buf2), .Y(_2710_) );
OAI21X1 OAI21X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_1617_), .B(raddr1_0_bF_buf9_), .C(raddr1_1_bF_buf10_bF_buf0_), .Y(_2711_) );
AOI21X1 AOI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(regs_16__6_), .B(raddr1_0_bF_buf8_), .C(_2711_), .Y(_2712_) );
NOR2X1 NOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf7_), .B(_1519_), .Y(_2713_) );
NAND2X1 NAND2X1_373 ( .gnd(gnd), .vdd(vdd), .A(regs_18__6_), .B(raddr1_0_bF_buf6_), .Y(_2714_) );
NAND2X1 NAND2X1_374 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf1), .B(_2714_), .Y(_2715_) );
OAI21X1 OAI21X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_2715_), .B(_2713_), .C(raddr1_2_bF_buf7_), .Y(_2716_) );
OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_2712_), .B(_2716_), .C(_2710_), .D(_2707_), .Y(_2717_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(regs_29__6_), .Y(_2718_) );
NAND2X1 NAND2X1_375 ( .gnd(gnd), .vdd(vdd), .A(regs_28__6_), .B(raddr1_0_bF_buf5_), .Y(_2719_) );
OAI21X1 OAI21X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_2718_), .B(raddr1_0_bF_buf4_), .C(_2719_), .Y(_2720_) );
MUX2X1 MUX2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_2720_), .B(regs_30__6_), .S(raddr1_1_bF_buf9_bF_buf0_), .Y(_2721_) );
NAND2X1 NAND2X1_376 ( .gnd(gnd), .vdd(vdd), .A(regs_26__6_), .B(raddr1_0_bF_buf3_), .Y(_2722_) );
OAI21X1 OAI21X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .B(raddr1_0_bF_buf2_), .C(_2722_), .Y(_2723_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(regs_25__6_), .Y(_2724_) );
NAND2X1 NAND2X1_377 ( .gnd(gnd), .vdd(vdd), .A(regs_24__6_), .B(raddr1_0_bF_buf1_), .Y(_2725_) );
OAI21X1 OAI21X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_2724_), .B(raddr1_0_bF_buf0_), .C(_2725_), .Y(_2726_) );
MUX2X1 MUX2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_2726_), .B(_2723_), .S(raddr1_1_bF_buf8_), .Y(_2727_) );
MUX2X1 MUX2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_2727_), .B(_2721_), .S(raddr1_2_bF_buf6_), .Y(_2728_) );
MUX2X1 MUX2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_2728_), .B(_2717_), .S(_2398__bF_buf1), .Y(_2729_) );
NAND2X1 NAND2X1_378 ( .gnd(gnd), .vdd(vdd), .A(regs_6__6_), .B(raddr1_0_bF_buf96_), .Y(_2730_) );
OAI21X1 OAI21X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_2113_), .B(raddr1_0_bF_buf95_), .C(_2730_), .Y(_2731_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(regs_5__6_), .Y(_2732_) );
NAND2X1 NAND2X1_379 ( .gnd(gnd), .vdd(vdd), .A(regs_4__6_), .B(raddr1_0_bF_buf94_), .Y(_2733_) );
OAI21X1 OAI21X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_2732_), .B(raddr1_0_bF_buf93_), .C(_2733_), .Y(_2734_) );
MUX2X1 MUX2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_2734_), .B(_2731_), .S(raddr1_1_bF_buf7_), .Y(_2735_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(regs_3__6_), .Y(_2736_) );
NAND2X1 NAND2X1_380 ( .gnd(gnd), .vdd(vdd), .A(regs_2__6_), .B(raddr1_0_bF_buf92_), .Y(_2737_) );
OAI21X1 OAI21X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_2736_), .B(raddr1_0_bF_buf91_), .C(_2737_), .Y(_2738_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(regs_1__6_), .Y(_2739_) );
NAND2X1 NAND2X1_381 ( .gnd(gnd), .vdd(vdd), .A(regs_0__6_), .B(raddr1_0_bF_buf90_), .Y(_2740_) );
OAI21X1 OAI21X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(raddr1_0_bF_buf89_), .C(_2740_), .Y(_2741_) );
MUX2X1 MUX2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_2741_), .B(_2738_), .S(raddr1_1_bF_buf6_), .Y(_2742_) );
MUX2X1 MUX2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_2742_), .B(_2735_), .S(raddr1_2_bF_buf5_), .Y(_2743_) );
NAND2X1 NAND2X1_382 ( .gnd(gnd), .vdd(vdd), .A(regs_14__6_), .B(raddr1_0_bF_buf88_), .Y(_2744_) );
OAI21X1 OAI21X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_1717_), .B(raddr1_0_bF_buf87_), .C(_2744_), .Y(_2745_) );
NAND2X1 NAND2X1_383 ( .gnd(gnd), .vdd(vdd), .A(regs_12__6_), .B(raddr1_0_bF_buf86_), .Y(_2746_) );
OAI21X1 OAI21X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_1815_), .B(raddr1_0_bF_buf85_), .C(_2746_), .Y(_2747_) );
MUX2X1 MUX2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_2747_), .B(_2745_), .S(raddr1_1_bF_buf5_), .Y(_2748_) );
NAND2X1 NAND2X1_384 ( .gnd(gnd), .vdd(vdd), .A(regs_10__6_), .B(raddr1_0_bF_buf84_), .Y(_2749_) );
OAI21X1 OAI21X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_1914_), .B(raddr1_0_bF_buf83_), .C(_2749_), .Y(_2750_) );
NAND2X1 NAND2X1_385 ( .gnd(gnd), .vdd(vdd), .A(regs_8__6_), .B(raddr1_0_bF_buf82_), .Y(_2751_) );
OAI21X1 OAI21X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_2012_), .B(raddr1_0_bF_buf81_), .C(_2751_), .Y(_2752_) );
MUX2X1 MUX2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_2752_), .B(_2750_), .S(raddr1_1_bF_buf4_), .Y(_2753_) );
MUX2X1 MUX2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_2753_), .B(_2748_), .S(raddr1_2_bF_buf4_), .Y(_2754_) );
MUX2X1 MUX2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_2754_), .B(_2743_), .S(_2398__bF_buf0), .Y(_2755_) );
MUX2X1 MUX2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_2755_), .B(_2729_), .S(raddr1_4_bF_buf3_), .Y(_5511__6_) );
NAND2X1 NAND2X1_386 ( .gnd(gnd), .vdd(vdd), .A(regs_22__7_), .B(raddr1_0_bF_buf80_), .Y(_2756_) );
OAI21X1 OAI21X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_1324_), .B(raddr1_0_bF_buf79_), .C(_2756_), .Y(_2757_) );
NAND2X1 NAND2X1_387 ( .gnd(gnd), .vdd(vdd), .A(regs_20__7_), .B(raddr1_0_bF_buf78_), .Y(_2758_) );
OAI21X1 OAI21X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_1422_), .B(raddr1_0_bF_buf77_), .C(_2758_), .Y(_2759_) );
MUX2X1 MUX2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_2759_), .B(_2757_), .S(raddr1_1_bF_buf3_), .Y(_2760_) );
NAND2X1 NAND2X1_388 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf1), .B(_2760_), .Y(_2761_) );
NAND2X1 NAND2X1_389 ( .gnd(gnd), .vdd(vdd), .A(regs_18__7_), .B(raddr1_0_bF_buf76_), .Y(_2762_) );
OAI21X1 OAI21X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_1521_), .B(raddr1_0_bF_buf75_), .C(_2762_), .Y(_2763_) );
NAND2X1 NAND2X1_390 ( .gnd(gnd), .vdd(vdd), .A(regs_16__7_), .B(raddr1_0_bF_buf74_), .Y(_2764_) );
OAI21X1 OAI21X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_1619_), .B(raddr1_0_bF_buf73_), .C(_2764_), .Y(_2765_) );
MUX2X1 MUX2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_2765_), .B(_2763_), .S(raddr1_1_bF_buf2_), .Y(_2766_) );
AOI21X1 AOI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(raddr1_2_bF_buf3_), .B(_2766_), .C(_2398__bF_buf7), .Y(_2767_) );
OAI21X1 OAI21X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_1157_), .B(raddr1_0_bF_buf72_), .C(raddr1_2_bF_buf2_), .Y(_2768_) );
AOI21X1 AOI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(regs_26__7_), .B(raddr1_0_bF_buf71_), .C(_2768_), .Y(_2769_) );
OAI21X1 OAI21X1_1169 ( .gnd(gnd), .vdd(vdd), .A(regs_30__7_), .B(raddr1_2_bF_buf1_), .C(_2415__bF_buf0), .Y(_2770_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(regs_25__7_), .Y(_2771_) );
OAI21X1 OAI21X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_2771_), .B(raddr1_0_bF_buf70_), .C(raddr1_2_bF_buf0_), .Y(_2772_) );
AOI21X1 AOI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(regs_24__7_), .B(raddr1_0_bF_buf69_), .C(_2772_), .Y(_2773_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(regs_29__7_), .Y(_2774_) );
NOR2X1 NOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf68_), .B(_2774_), .Y(_2775_) );
NAND2X1 NAND2X1_391 ( .gnd(gnd), .vdd(vdd), .A(regs_28__7_), .B(raddr1_0_bF_buf67_), .Y(_2776_) );
NAND2X1 NAND2X1_392 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf0), .B(_2776_), .Y(_2777_) );
OAI21X1 OAI21X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_2777_), .B(_2775_), .C(raddr1_1_bF_buf1_), .Y(_2778_) );
OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_2769_), .B(_2770_), .C(_2778_), .D(_2773_), .Y(_2779_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_2779_), .B(_2398__bF_buf6), .C(_2761_), .D(_2767_), .Y(_2780_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(regs_5__7_), .Y(_2781_) );
OAI21X1 OAI21X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_2781_), .B(raddr1_0_bF_buf66_), .C(raddr1_1_bF_buf0_), .Y(_2782_) );
AOI21X1 AOI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(regs_4__7_), .B(raddr1_0_bF_buf65_), .C(_2782_), .Y(_2783_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(regs_6__7_), .B(raddr1_0_bF_buf64_), .Y(_2784_) );
OAI21X1 OAI21X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_2115_), .B(raddr1_0_bF_buf63_), .C(_2415__bF_buf8), .Y(_2785_) );
OAI21X1 OAI21X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_2785_), .B(_2784_), .C(_2399__bF_buf8), .Y(_2786_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(regs_1__7_), .Y(_2787_) );
OAI21X1 OAI21X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_2787_), .B(raddr1_0_bF_buf62_), .C(raddr1_1_bF_buf14_bF_buf3_), .Y(_2788_) );
AOI21X1 AOI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(regs_0__7_), .B(raddr1_0_bF_buf61_), .C(_2788_), .Y(_2789_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(regs_3__7_), .Y(_2790_) );
NOR2X1 NOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf60_), .B(_2790_), .Y(_2791_) );
NAND2X1 NAND2X1_393 ( .gnd(gnd), .vdd(vdd), .A(regs_2__7_), .B(raddr1_0_bF_buf59_), .Y(_2792_) );
NAND2X1 NAND2X1_394 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf7), .B(_2792_), .Y(_2793_) );
OAI21X1 OAI21X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_2793_), .B(_2791_), .C(raddr1_2_bF_buf10_), .Y(_2794_) );
OAI22X1 OAI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_2789_), .B(_2794_), .C(_2786_), .D(_2783_), .Y(_2795_) );
NAND2X1 NAND2X1_395 ( .gnd(gnd), .vdd(vdd), .A(regs_10__7_), .B(raddr1_0_bF_buf58_), .Y(_2796_) );
OAI21X1 OAI21X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_1916_), .B(raddr1_0_bF_buf57_), .C(_2796_), .Y(_2797_) );
NAND2X1 NAND2X1_396 ( .gnd(gnd), .vdd(vdd), .A(regs_8__7_), .B(raddr1_0_bF_buf56_), .Y(_2798_) );
OAI21X1 OAI21X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_2014_), .B(raddr1_0_bF_buf55_), .C(_2798_), .Y(_2799_) );
MUX2X1 MUX2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_2799_), .B(_2797_), .S(raddr1_1_bF_buf13_bF_buf3_), .Y(_2800_) );
NAND2X1 NAND2X1_397 ( .gnd(gnd), .vdd(vdd), .A(regs_14__7_), .B(raddr1_0_bF_buf54_), .Y(_2801_) );
OAI21X1 OAI21X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_1719_), .B(raddr1_0_bF_buf53_), .C(_2801_), .Y(_2802_) );
NAND2X1 NAND2X1_398 ( .gnd(gnd), .vdd(vdd), .A(regs_12__7_), .B(raddr1_0_bF_buf52_), .Y(_2803_) );
OAI21X1 OAI21X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_1817_), .B(raddr1_0_bF_buf51_), .C(_2803_), .Y(_2804_) );
MUX2X1 MUX2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_2804_), .B(_2802_), .S(raddr1_1_bF_buf12_bF_buf3_), .Y(_2805_) );
MUX2X1 MUX2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_2805_), .B(_2800_), .S(_2399__bF_buf7), .Y(_2806_) );
MUX2X1 MUX2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_2806_), .B(_2795_), .S(_2398__bF_buf5), .Y(_2807_) );
MUX2X1 MUX2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_2807_), .B(_2780_), .S(raddr1_4_bF_buf2_), .Y(_5511__7_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(regs_5__8_), .Y(_2808_) );
OAI21X1 OAI21X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_2808_), .B(raddr1_0_bF_buf50_), .C(raddr1_1_bF_buf11_bF_buf3_), .Y(_2809_) );
AOI21X1 AOI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(regs_4__8_), .B(raddr1_0_bF_buf49_), .C(_2809_), .Y(_2810_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(regs_6__8_), .B(raddr1_0_bF_buf48_), .Y(_2811_) );
OAI21X1 OAI21X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_2117_), .B(raddr1_0_bF_buf47_), .C(_2415__bF_buf6), .Y(_2812_) );
OAI21X1 OAI21X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_2812_), .B(_2811_), .C(_2399__bF_buf6), .Y(_2813_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(regs_1__8_), .Y(_2814_) );
OAI21X1 OAI21X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_2814_), .B(raddr1_0_bF_buf46_), .C(raddr1_1_bF_buf10_bF_buf3_), .Y(_2815_) );
AOI21X1 AOI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(regs_0__8_), .B(raddr1_0_bF_buf45_), .C(_2815_), .Y(_2816_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(regs_3__8_), .Y(_2817_) );
NOR2X1 NOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf44_), .B(_2817_), .Y(_2818_) );
NAND2X1 NAND2X1_399 ( .gnd(gnd), .vdd(vdd), .A(regs_2__8_), .B(raddr1_0_bF_buf43_), .Y(_2819_) );
NAND2X1 NAND2X1_400 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf5), .B(_2819_), .Y(_2820_) );
OAI21X1 OAI21X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_2820_), .B(_2818_), .C(raddr1_2_bF_buf9_), .Y(_2821_) );
OAI22X1 OAI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_2816_), .B(_2821_), .C(_2813_), .D(_2810_), .Y(_2822_) );
NAND2X1 NAND2X1_401 ( .gnd(gnd), .vdd(vdd), .A(regs_10__8_), .B(raddr1_0_bF_buf42_), .Y(_2823_) );
OAI21X1 OAI21X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_1918_), .B(raddr1_0_bF_buf41_), .C(_2823_), .Y(_2824_) );
NAND2X1 NAND2X1_402 ( .gnd(gnd), .vdd(vdd), .A(regs_8__8_), .B(raddr1_0_bF_buf40_), .Y(_2825_) );
OAI21X1 OAI21X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_2016_), .B(raddr1_0_bF_buf39_), .C(_2825_), .Y(_2826_) );
MUX2X1 MUX2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_2826_), .B(_2824_), .S(raddr1_1_bF_buf9_bF_buf3_), .Y(_2827_) );
NAND2X1 NAND2X1_403 ( .gnd(gnd), .vdd(vdd), .A(regs_14__8_), .B(raddr1_0_bF_buf38_), .Y(_2828_) );
OAI21X1 OAI21X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_1721_), .B(raddr1_0_bF_buf37_), .C(_2828_), .Y(_2829_) );
NAND2X1 NAND2X1_404 ( .gnd(gnd), .vdd(vdd), .A(regs_12__8_), .B(raddr1_0_bF_buf36_), .Y(_2830_) );
OAI21X1 OAI21X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_1819_), .B(raddr1_0_bF_buf35_), .C(_2830_), .Y(_2831_) );
MUX2X1 MUX2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_2831_), .B(_2829_), .S(raddr1_1_bF_buf8_), .Y(_2832_) );
MUX2X1 MUX2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_2832_), .B(_2827_), .S(_2399__bF_buf5), .Y(_2833_) );
MUX2X1 MUX2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_2833_), .B(_2822_), .S(_2398__bF_buf4), .Y(_2834_) );
OAI21X1 OAI21X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .B(raddr1_0_bF_buf34_), .C(raddr1_1_bF_buf7_), .Y(_2835_) );
AOI21X1 AOI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(regs_16__8_), .B(raddr1_0_bF_buf33_), .C(_2835_), .Y(_2836_) );
NOR2X1 NOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf32_), .B(_1523_), .Y(_2837_) );
NAND2X1 NAND2X1_405 ( .gnd(gnd), .vdd(vdd), .A(regs_18__8_), .B(raddr1_0_bF_buf31_), .Y(_2838_) );
NAND2X1 NAND2X1_406 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf4), .B(_2838_), .Y(_2839_) );
OAI21X1 OAI21X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_2839_), .B(_2837_), .C(raddr1_2_bF_buf8_), .Y(_2840_) );
OAI21X1 OAI21X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_1424_), .B(raddr1_0_bF_buf30_), .C(raddr1_1_bF_buf6_), .Y(_2841_) );
AOI21X1 AOI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(regs_20__8_), .B(raddr1_0_bF_buf29_), .C(_2841_), .Y(_2842_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(regs_22__8_), .B(raddr1_0_bF_buf28_), .Y(_2843_) );
OAI21X1 OAI21X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_1326_), .B(raddr1_0_bF_buf27_), .C(_2415__bF_buf3), .Y(_2844_) );
OAI21X1 OAI21X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_2844_), .B(_2843_), .C(_2399__bF_buf4), .Y(_2845_) );
OAI22X1 OAI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_2836_), .B(_2840_), .C(_2845_), .D(_2842_), .Y(_2846_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(regs_29__8_), .Y(_2847_) );
NAND2X1 NAND2X1_407 ( .gnd(gnd), .vdd(vdd), .A(regs_28__8_), .B(raddr1_0_bF_buf26_), .Y(_2848_) );
OAI21X1 OAI21X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_2847_), .B(raddr1_0_bF_buf25_), .C(_2848_), .Y(_2849_) );
MUX2X1 MUX2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_2849_), .B(regs_30__8_), .S(raddr1_1_bF_buf5_), .Y(_2850_) );
NAND2X1 NAND2X1_408 ( .gnd(gnd), .vdd(vdd), .A(regs_26__8_), .B(raddr1_0_bF_buf24_), .Y(_2851_) );
OAI21X1 OAI21X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_1159_), .B(raddr1_0_bF_buf23_), .C(_2851_), .Y(_2852_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(regs_25__8_), .Y(_2853_) );
NAND2X1 NAND2X1_409 ( .gnd(gnd), .vdd(vdd), .A(regs_24__8_), .B(raddr1_0_bF_buf22_), .Y(_2854_) );
OAI21X1 OAI21X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_2853_), .B(raddr1_0_bF_buf21_), .C(_2854_), .Y(_2855_) );
MUX2X1 MUX2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_2855_), .B(_2852_), .S(raddr1_1_bF_buf4_), .Y(_2856_) );
MUX2X1 MUX2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_2856_), .B(_2850_), .S(raddr1_2_bF_buf7_), .Y(_2857_) );
MUX2X1 MUX2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_2857_), .B(_2846_), .S(_2398__bF_buf3), .Y(_2858_) );
MUX2X1 MUX2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_2834_), .B(_2858_), .S(raddr1_4_bF_buf1_), .Y(_5511__8_) );
NAND2X1 NAND2X1_410 ( .gnd(gnd), .vdd(vdd), .A(regs_22__9_), .B(raddr1_0_bF_buf20_), .Y(_2859_) );
OAI21X1 OAI21X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_1328_), .B(raddr1_0_bF_buf19_), .C(_2859_), .Y(_2860_) );
NAND2X1 NAND2X1_411 ( .gnd(gnd), .vdd(vdd), .A(regs_20__9_), .B(raddr1_0_bF_buf18_), .Y(_2861_) );
OAI21X1 OAI21X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_1426_), .B(raddr1_0_bF_buf17_), .C(_2861_), .Y(_2862_) );
MUX2X1 MUX2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_2862_), .B(_2860_), .S(raddr1_1_bF_buf3_), .Y(_2863_) );
NAND2X1 NAND2X1_412 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf3), .B(_2863_), .Y(_2864_) );
NAND2X1 NAND2X1_413 ( .gnd(gnd), .vdd(vdd), .A(regs_18__9_), .B(raddr1_0_bF_buf16_), .Y(_2865_) );
OAI21X1 OAI21X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_1525_), .B(raddr1_0_bF_buf15_), .C(_2865_), .Y(_2866_) );
NAND2X1 NAND2X1_414 ( .gnd(gnd), .vdd(vdd), .A(regs_16__9_), .B(raddr1_0_bF_buf14_), .Y(_2867_) );
OAI21X1 OAI21X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(raddr1_0_bF_buf13_), .C(_2867_), .Y(_2868_) );
MUX2X1 MUX2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_2868_), .B(_2866_), .S(raddr1_1_bF_buf2_), .Y(_2869_) );
AOI21X1 AOI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(raddr1_2_bF_buf6_), .B(_2869_), .C(_2398__bF_buf2), .Y(_2870_) );
OAI21X1 OAI21X1_1202 ( .gnd(gnd), .vdd(vdd), .A(_1161_), .B(raddr1_0_bF_buf12_), .C(raddr1_2_bF_buf5_), .Y(_2871_) );
AOI21X1 AOI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(regs_26__9_), .B(raddr1_0_bF_buf11_), .C(_2871_), .Y(_2872_) );
OAI21X1 OAI21X1_1203 ( .gnd(gnd), .vdd(vdd), .A(regs_30__9_), .B(raddr1_2_bF_buf4_), .C(_2415__bF_buf2), .Y(_2873_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(regs_25__9_), .Y(_2874_) );
OAI21X1 OAI21X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_2874_), .B(raddr1_0_bF_buf10_), .C(raddr1_2_bF_buf3_), .Y(_2875_) );
AOI21X1 AOI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(regs_24__9_), .B(raddr1_0_bF_buf9_), .C(_2875_), .Y(_2876_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(regs_29__9_), .Y(_2877_) );
NOR2X1 NOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf8_), .B(_2877_), .Y(_2878_) );
NAND2X1 NAND2X1_415 ( .gnd(gnd), .vdd(vdd), .A(regs_28__9_), .B(raddr1_0_bF_buf7_), .Y(_2879_) );
NAND2X1 NAND2X1_416 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf2), .B(_2879_), .Y(_2880_) );
OAI21X1 OAI21X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_2880_), .B(_2878_), .C(raddr1_1_bF_buf1_), .Y(_2881_) );
OAI22X1 OAI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_2872_), .B(_2873_), .C(_2881_), .D(_2876_), .Y(_2882_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_2882_), .B(_2398__bF_buf1), .C(_2864_), .D(_2870_), .Y(_2883_) );
NAND2X1 NAND2X1_417 ( .gnd(gnd), .vdd(vdd), .A(regs_6__9_), .B(raddr1_0_bF_buf6_), .Y(_2884_) );
OAI21X1 OAI21X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_2119_), .B(raddr1_0_bF_buf5_), .C(_2884_), .Y(_2885_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(regs_5__9_), .Y(_2886_) );
NAND2X1 NAND2X1_418 ( .gnd(gnd), .vdd(vdd), .A(regs_4__9_), .B(raddr1_0_bF_buf4_), .Y(_2887_) );
OAI21X1 OAI21X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_2886_), .B(raddr1_0_bF_buf3_), .C(_2887_), .Y(_2888_) );
MUX2X1 MUX2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_2888_), .B(_2885_), .S(raddr1_1_bF_buf0_), .Y(_2889_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(regs_3__9_), .Y(_2890_) );
NAND2X1 NAND2X1_419 ( .gnd(gnd), .vdd(vdd), .A(regs_2__9_), .B(raddr1_0_bF_buf2_), .Y(_2891_) );
OAI21X1 OAI21X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_2890_), .B(raddr1_0_bF_buf1_), .C(_2891_), .Y(_2892_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(regs_1__9_), .Y(_2893_) );
NAND2X1 NAND2X1_420 ( .gnd(gnd), .vdd(vdd), .A(regs_0__9_), .B(raddr1_0_bF_buf0_), .Y(_2894_) );
OAI21X1 OAI21X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_2893_), .B(raddr1_0_bF_buf96_), .C(_2894_), .Y(_2895_) );
MUX2X1 MUX2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_2895_), .B(_2892_), .S(raddr1_1_bF_buf14_bF_buf2_), .Y(_2896_) );
MUX2X1 MUX2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_2896_), .B(_2889_), .S(raddr1_2_bF_buf2_), .Y(_2897_) );
NAND2X1 NAND2X1_421 ( .gnd(gnd), .vdd(vdd), .A(regs_14__9_), .B(raddr1_0_bF_buf95_), .Y(_2898_) );
OAI21X1 OAI21X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_1723_), .B(raddr1_0_bF_buf94_), .C(_2898_), .Y(_2899_) );
NAND2X1 NAND2X1_422 ( .gnd(gnd), .vdd(vdd), .A(regs_12__9_), .B(raddr1_0_bF_buf93_), .Y(_2900_) );
OAI21X1 OAI21X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_1821_), .B(raddr1_0_bF_buf92_), .C(_2900_), .Y(_2901_) );
MUX2X1 MUX2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_2901_), .B(_2899_), .S(raddr1_1_bF_buf13_bF_buf2_), .Y(_2902_) );
NAND2X1 NAND2X1_423 ( .gnd(gnd), .vdd(vdd), .A(regs_10__9_), .B(raddr1_0_bF_buf91_), .Y(_2903_) );
OAI21X1 OAI21X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_1920_), .B(raddr1_0_bF_buf90_), .C(_2903_), .Y(_2904_) );
NAND2X1 NAND2X1_424 ( .gnd(gnd), .vdd(vdd), .A(regs_8__9_), .B(raddr1_0_bF_buf89_), .Y(_2905_) );
OAI21X1 OAI21X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_2018_), .B(raddr1_0_bF_buf88_), .C(_2905_), .Y(_2906_) );
MUX2X1 MUX2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_2906_), .B(_2904_), .S(raddr1_1_bF_buf12_bF_buf2_), .Y(_2907_) );
MUX2X1 MUX2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_2907_), .B(_2902_), .S(raddr1_2_bF_buf1_), .Y(_2908_) );
MUX2X1 MUX2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_2908_), .B(_2897_), .S(_2398__bF_buf0), .Y(_2909_) );
MUX2X1 MUX2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_2909_), .B(_2883_), .S(raddr1_4_bF_buf0_), .Y(_5511__9_) );
NAND2X1 NAND2X1_425 ( .gnd(gnd), .vdd(vdd), .A(regs_22__10_), .B(raddr1_0_bF_buf87_), .Y(_2910_) );
OAI21X1 OAI21X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_1330_), .B(raddr1_0_bF_buf86_), .C(_2910_), .Y(_2911_) );
NAND2X1 NAND2X1_426 ( .gnd(gnd), .vdd(vdd), .A(regs_20__10_), .B(raddr1_0_bF_buf85_), .Y(_2912_) );
OAI21X1 OAI21X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_1428_), .B(raddr1_0_bF_buf84_), .C(_2912_), .Y(_2913_) );
MUX2X1 MUX2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_2913_), .B(_2911_), .S(raddr1_1_bF_buf11_bF_buf2_), .Y(_2914_) );
NAND2X1 NAND2X1_427 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf1), .B(_2914_), .Y(_2915_) );
NAND2X1 NAND2X1_428 ( .gnd(gnd), .vdd(vdd), .A(regs_18__10_), .B(raddr1_0_bF_buf83_), .Y(_2916_) );
OAI21X1 OAI21X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_1527_), .B(raddr1_0_bF_buf82_), .C(_2916_), .Y(_2917_) );
NAND2X1 NAND2X1_429 ( .gnd(gnd), .vdd(vdd), .A(regs_16__10_), .B(raddr1_0_bF_buf81_), .Y(_2918_) );
OAI21X1 OAI21X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_1625_), .B(raddr1_0_bF_buf80_), .C(_2918_), .Y(_2919_) );
MUX2X1 MUX2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_2919_), .B(_2917_), .S(raddr1_1_bF_buf10_bF_buf2_), .Y(_2920_) );
AOI21X1 AOI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(raddr1_2_bF_buf0_), .B(_2920_), .C(_2398__bF_buf7), .Y(_2921_) );
OAI21X1 OAI21X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(raddr1_0_bF_buf79_), .C(raddr1_2_bF_buf10_), .Y(_2922_) );
AOI21X1 AOI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(regs_26__10_), .B(raddr1_0_bF_buf78_), .C(_2922_), .Y(_2923_) );
OAI21X1 OAI21X1_1219 ( .gnd(gnd), .vdd(vdd), .A(regs_30__10_), .B(raddr1_2_bF_buf9_), .C(_2415__bF_buf1), .Y(_2924_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(regs_25__10_), .Y(_2925_) );
OAI21X1 OAI21X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_2925_), .B(raddr1_0_bF_buf77_), .C(raddr1_2_bF_buf8_), .Y(_2926_) );
AOI21X1 AOI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(regs_24__10_), .B(raddr1_0_bF_buf76_), .C(_2926_), .Y(_2927_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(regs_29__10_), .Y(_2928_) );
NOR2X1 NOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf75_), .B(_2928_), .Y(_2929_) );
NAND2X1 NAND2X1_430 ( .gnd(gnd), .vdd(vdd), .A(regs_28__10_), .B(raddr1_0_bF_buf74_), .Y(_2930_) );
NAND2X1 NAND2X1_431 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf0), .B(_2930_), .Y(_2931_) );
OAI21X1 OAI21X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_2931_), .B(_2929_), .C(raddr1_1_bF_buf9_bF_buf2_), .Y(_2932_) );
OAI22X1 OAI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_2923_), .B(_2924_), .C(_2932_), .D(_2927_), .Y(_2933_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_2933_), .B(_2398__bF_buf6), .C(_2915_), .D(_2921_), .Y(_2934_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(regs_5__10_), .Y(_2935_) );
OAI21X1 OAI21X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_2935_), .B(raddr1_0_bF_buf73_), .C(raddr1_1_bF_buf8_), .Y(_2936_) );
AOI21X1 AOI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(regs_4__10_), .B(raddr1_0_bF_buf72_), .C(_2936_), .Y(_2937_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(regs_6__10_), .B(raddr1_0_bF_buf71_), .Y(_2938_) );
OAI21X1 OAI21X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_2121_), .B(raddr1_0_bF_buf70_), .C(_2415__bF_buf0), .Y(_2939_) );
OAI21X1 OAI21X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_2939_), .B(_2938_), .C(_2399__bF_buf8), .Y(_2940_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(regs_1__10_), .Y(_2941_) );
OAI21X1 OAI21X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_2941_), .B(raddr1_0_bF_buf69_), .C(raddr1_1_bF_buf7_), .Y(_2942_) );
AOI21X1 AOI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(regs_0__10_), .B(raddr1_0_bF_buf68_), .C(_2942_), .Y(_2943_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(regs_3__10_), .Y(_2944_) );
NOR2X1 NOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf67_), .B(_2944_), .Y(_2945_) );
NAND2X1 NAND2X1_432 ( .gnd(gnd), .vdd(vdd), .A(regs_2__10_), .B(raddr1_0_bF_buf66_), .Y(_2946_) );
NAND2X1 NAND2X1_433 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf8), .B(_2946_), .Y(_2947_) );
OAI21X1 OAI21X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_2947_), .B(_2945_), .C(raddr1_2_bF_buf7_), .Y(_2948_) );
OAI22X1 OAI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_2943_), .B(_2948_), .C(_2940_), .D(_2937_), .Y(_2949_) );
NAND2X1 NAND2X1_434 ( .gnd(gnd), .vdd(vdd), .A(regs_10__10_), .B(raddr1_0_bF_buf65_), .Y(_2950_) );
OAI21X1 OAI21X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_1922_), .B(raddr1_0_bF_buf64_), .C(_2950_), .Y(_2951_) );
NAND2X1 NAND2X1_435 ( .gnd(gnd), .vdd(vdd), .A(regs_8__10_), .B(raddr1_0_bF_buf63_), .Y(_2952_) );
OAI21X1 OAI21X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_2020_), .B(raddr1_0_bF_buf62_), .C(_2952_), .Y(_2953_) );
MUX2X1 MUX2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_2953_), .B(_2951_), .S(raddr1_1_bF_buf6_), .Y(_2954_) );
NAND2X1 NAND2X1_436 ( .gnd(gnd), .vdd(vdd), .A(regs_14__10_), .B(raddr1_0_bF_buf61_), .Y(_2955_) );
OAI21X1 OAI21X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_1725_), .B(raddr1_0_bF_buf60_), .C(_2955_), .Y(_2956_) );
NAND2X1 NAND2X1_437 ( .gnd(gnd), .vdd(vdd), .A(regs_12__10_), .B(raddr1_0_bF_buf59_), .Y(_2957_) );
OAI21X1 OAI21X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_1823_), .B(raddr1_0_bF_buf58_), .C(_2957_), .Y(_2958_) );
MUX2X1 MUX2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_2958_), .B(_2956_), .S(raddr1_1_bF_buf5_), .Y(_2959_) );
MUX2X1 MUX2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_2959_), .B(_2954_), .S(_2399__bF_buf7), .Y(_2960_) );
MUX2X1 MUX2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_2960_), .B(_2949_), .S(_2398__bF_buf5), .Y(_2961_) );
MUX2X1 MUX2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_2961_), .B(_2934_), .S(raddr1_4_bF_buf4_), .Y(_5511__10_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(regs_5__11_), .Y(_2962_) );
OAI21X1 OAI21X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_2962_), .B(raddr1_0_bF_buf57_), .C(raddr1_1_bF_buf4_), .Y(_2963_) );
AOI21X1 AOI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(regs_4__11_), .B(raddr1_0_bF_buf56_), .C(_2963_), .Y(_2964_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(regs_6__11_), .B(raddr1_0_bF_buf55_), .Y(_2965_) );
OAI21X1 OAI21X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_2123_), .B(raddr1_0_bF_buf54_), .C(_2415__bF_buf7), .Y(_2966_) );
OAI21X1 OAI21X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_2966_), .B(_2965_), .C(_2399__bF_buf6), .Y(_2967_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(regs_1__11_), .Y(_2968_) );
OAI21X1 OAI21X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_2968_), .B(raddr1_0_bF_buf53_), .C(raddr1_1_bF_buf3_), .Y(_2969_) );
AOI21X1 AOI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(regs_0__11_), .B(raddr1_0_bF_buf52_), .C(_2969_), .Y(_2970_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(regs_3__11_), .Y(_2971_) );
NOR2X1 NOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf51_), .B(_2971_), .Y(_2972_) );
NAND2X1 NAND2X1_438 ( .gnd(gnd), .vdd(vdd), .A(regs_2__11_), .B(raddr1_0_bF_buf50_), .Y(_2973_) );
NAND2X1 NAND2X1_439 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf6), .B(_2973_), .Y(_2974_) );
OAI21X1 OAI21X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_2974_), .B(_2972_), .C(raddr1_2_bF_buf6_), .Y(_2975_) );
OAI22X1 OAI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_2970_), .B(_2975_), .C(_2967_), .D(_2964_), .Y(_2976_) );
NAND2X1 NAND2X1_440 ( .gnd(gnd), .vdd(vdd), .A(regs_10__11_), .B(raddr1_0_bF_buf49_), .Y(_2977_) );
OAI21X1 OAI21X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_1924_), .B(raddr1_0_bF_buf48_), .C(_2977_), .Y(_2978_) );
NAND2X1 NAND2X1_441 ( .gnd(gnd), .vdd(vdd), .A(regs_8__11_), .B(raddr1_0_bF_buf47_), .Y(_2979_) );
OAI21X1 OAI21X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_2022_), .B(raddr1_0_bF_buf46_), .C(_2979_), .Y(_2980_) );
MUX2X1 MUX2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_2980_), .B(_2978_), .S(raddr1_1_bF_buf2_), .Y(_2981_) );
NAND2X1 NAND2X1_442 ( .gnd(gnd), .vdd(vdd), .A(regs_14__11_), .B(raddr1_0_bF_buf45_), .Y(_2982_) );
OAI21X1 OAI21X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_1727_), .B(raddr1_0_bF_buf44_), .C(_2982_), .Y(_2983_) );
NAND2X1 NAND2X1_443 ( .gnd(gnd), .vdd(vdd), .A(regs_12__11_), .B(raddr1_0_bF_buf43_), .Y(_2984_) );
OAI21X1 OAI21X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_1825_), .B(raddr1_0_bF_buf42_), .C(_2984_), .Y(_2985_) );
MUX2X1 MUX2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_2985_), .B(_2983_), .S(raddr1_1_bF_buf1_), .Y(_2986_) );
MUX2X1 MUX2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_2986_), .B(_2981_), .S(_2399__bF_buf5), .Y(_2987_) );
MUX2X1 MUX2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_2987_), .B(_2976_), .S(_2398__bF_buf4), .Y(_2988_) );
OAI21X1 OAI21X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_1627_), .B(raddr1_0_bF_buf41_), .C(raddr1_1_bF_buf0_), .Y(_2989_) );
AOI21X1 AOI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(regs_16__11_), .B(raddr1_0_bF_buf40_), .C(_2989_), .Y(_2990_) );
NOR2X1 NOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf39_), .B(_1529_), .Y(_2991_) );
NAND2X1 NAND2X1_444 ( .gnd(gnd), .vdd(vdd), .A(regs_18__11_), .B(raddr1_0_bF_buf38_), .Y(_2992_) );
NAND2X1 NAND2X1_445 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf5), .B(_2992_), .Y(_2993_) );
OAI21X1 OAI21X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_2993_), .B(_2991_), .C(raddr1_2_bF_buf5_), .Y(_2994_) );
OAI21X1 OAI21X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_1430_), .B(raddr1_0_bF_buf37_), .C(raddr1_1_bF_buf14_bF_buf1_), .Y(_2995_) );
AOI21X1 AOI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(regs_20__11_), .B(raddr1_0_bF_buf36_), .C(_2995_), .Y(_2996_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(regs_22__11_), .B(raddr1_0_bF_buf35_), .Y(_2997_) );
OAI21X1 OAI21X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_1332_), .B(raddr1_0_bF_buf34_), .C(_2415__bF_buf4), .Y(_2998_) );
OAI21X1 OAI21X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_2998_), .B(_2997_), .C(_2399__bF_buf4), .Y(_2999_) );
OAI22X1 OAI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_2990_), .B(_2994_), .C(_2999_), .D(_2996_), .Y(_3000_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(regs_29__11_), .Y(_3001_) );
NAND2X1 NAND2X1_446 ( .gnd(gnd), .vdd(vdd), .A(regs_28__11_), .B(raddr1_0_bF_buf33_), .Y(_3002_) );
OAI21X1 OAI21X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_3001_), .B(raddr1_0_bF_buf32_), .C(_3002_), .Y(_3003_) );
MUX2X1 MUX2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_3003_), .B(regs_30__11_), .S(raddr1_1_bF_buf13_bF_buf1_), .Y(_3004_) );
NAND2X1 NAND2X1_447 ( .gnd(gnd), .vdd(vdd), .A(regs_26__11_), .B(raddr1_0_bF_buf31_), .Y(_3005_) );
OAI21X1 OAI21X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_1165_), .B(raddr1_0_bF_buf30_), .C(_3005_), .Y(_3006_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(regs_25__11_), .Y(_3007_) );
NAND2X1 NAND2X1_448 ( .gnd(gnd), .vdd(vdd), .A(regs_24__11_), .B(raddr1_0_bF_buf29_), .Y(_3008_) );
OAI21X1 OAI21X1_1247 ( .gnd(gnd), .vdd(vdd), .A(_3007_), .B(raddr1_0_bF_buf28_), .C(_3008_), .Y(_3009_) );
MUX2X1 MUX2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_3009_), .B(_3006_), .S(raddr1_1_bF_buf12_bF_buf1_), .Y(_3010_) );
MUX2X1 MUX2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_3010_), .B(_3004_), .S(raddr1_2_bF_buf4_), .Y(_3011_) );
MUX2X1 MUX2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_3011_), .B(_3000_), .S(_2398__bF_buf3), .Y(_3012_) );
MUX2X1 MUX2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_2988_), .B(_3012_), .S(raddr1_4_bF_buf3_), .Y(_5511__11_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(regs_5__12_), .Y(_3013_) );
OAI21X1 OAI21X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_3013_), .B(raddr1_0_bF_buf27_), .C(raddr1_1_bF_buf11_bF_buf1_), .Y(_3014_) );
AOI21X1 AOI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(regs_4__12_), .B(raddr1_0_bF_buf26_), .C(_3014_), .Y(_3015_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(regs_6__12_), .B(raddr1_0_bF_buf25_), .Y(_3016_) );
OAI21X1 OAI21X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_2125_), .B(raddr1_0_bF_buf24_), .C(_2415__bF_buf3), .Y(_3017_) );
OAI21X1 OAI21X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_3017_), .B(_3016_), .C(_2399__bF_buf3), .Y(_3018_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(regs_1__12_), .Y(_3019_) );
OAI21X1 OAI21X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_3019_), .B(raddr1_0_bF_buf23_), .C(raddr1_1_bF_buf10_bF_buf1_), .Y(_3020_) );
AOI21X1 AOI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(regs_0__12_), .B(raddr1_0_bF_buf22_), .C(_3020_), .Y(_3021_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(regs_3__12_), .Y(_3022_) );
NOR2X1 NOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf21_), .B(_3022_), .Y(_3023_) );
NAND2X1 NAND2X1_449 ( .gnd(gnd), .vdd(vdd), .A(regs_2__12_), .B(raddr1_0_bF_buf20_), .Y(_3024_) );
NAND2X1 NAND2X1_450 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf2), .B(_3024_), .Y(_3025_) );
OAI21X1 OAI21X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_3025_), .B(_3023_), .C(raddr1_2_bF_buf3_), .Y(_3026_) );
OAI22X1 OAI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_3021_), .B(_3026_), .C(_3018_), .D(_3015_), .Y(_3027_) );
NAND2X1 NAND2X1_451 ( .gnd(gnd), .vdd(vdd), .A(regs_10__12_), .B(raddr1_0_bF_buf19_), .Y(_3028_) );
OAI21X1 OAI21X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_1926_), .B(raddr1_0_bF_buf18_), .C(_3028_), .Y(_3029_) );
NAND2X1 NAND2X1_452 ( .gnd(gnd), .vdd(vdd), .A(regs_8__12_), .B(raddr1_0_bF_buf17_), .Y(_3030_) );
OAI21X1 OAI21X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_2024_), .B(raddr1_0_bF_buf16_), .C(_3030_), .Y(_3031_) );
MUX2X1 MUX2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_3031_), .B(_3029_), .S(raddr1_1_bF_buf9_bF_buf1_), .Y(_3032_) );
NAND2X1 NAND2X1_453 ( .gnd(gnd), .vdd(vdd), .A(regs_14__12_), .B(raddr1_0_bF_buf15_), .Y(_3033_) );
OAI21X1 OAI21X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_1729_), .B(raddr1_0_bF_buf14_), .C(_3033_), .Y(_3034_) );
NAND2X1 NAND2X1_454 ( .gnd(gnd), .vdd(vdd), .A(regs_12__12_), .B(raddr1_0_bF_buf13_), .Y(_3035_) );
OAI21X1 OAI21X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .B(raddr1_0_bF_buf12_), .C(_3035_), .Y(_3036_) );
MUX2X1 MUX2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_3036_), .B(_3034_), .S(raddr1_1_bF_buf8_), .Y(_3037_) );
MUX2X1 MUX2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_3037_), .B(_3032_), .S(_2399__bF_buf2), .Y(_3038_) );
MUX2X1 MUX2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_3038_), .B(_3027_), .S(_2398__bF_buf2), .Y(_3039_) );
OAI21X1 OAI21X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_1629_), .B(raddr1_0_bF_buf11_), .C(raddr1_1_bF_buf7_), .Y(_3040_) );
AOI21X1 AOI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(regs_16__12_), .B(raddr1_0_bF_buf10_), .C(_3040_), .Y(_3041_) );
NOR2X1 NOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf9_), .B(_1531_), .Y(_3042_) );
NAND2X1 NAND2X1_455 ( .gnd(gnd), .vdd(vdd), .A(regs_18__12_), .B(raddr1_0_bF_buf8_), .Y(_3043_) );
NAND2X1 NAND2X1_456 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf1), .B(_3043_), .Y(_3044_) );
OAI21X1 OAI21X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_3044_), .B(_3042_), .C(raddr1_2_bF_buf2_), .Y(_3045_) );
OAI21X1 OAI21X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_1432_), .B(raddr1_0_bF_buf7_), .C(raddr1_1_bF_buf6_), .Y(_3046_) );
AOI21X1 AOI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(regs_20__12_), .B(raddr1_0_bF_buf6_), .C(_3046_), .Y(_3047_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(regs_22__12_), .B(raddr1_0_bF_buf5_), .Y(_3048_) );
OAI21X1 OAI21X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_1334_), .B(raddr1_0_bF_buf4_), .C(_2415__bF_buf0), .Y(_3049_) );
OAI21X1 OAI21X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_3049_), .B(_3048_), .C(_2399__bF_buf1), .Y(_3050_) );
OAI22X1 OAI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_3041_), .B(_3045_), .C(_3050_), .D(_3047_), .Y(_3051_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(regs_29__12_), .Y(_3052_) );
NAND2X1 NAND2X1_457 ( .gnd(gnd), .vdd(vdd), .A(regs_28__12_), .B(raddr1_0_bF_buf3_), .Y(_3053_) );
OAI21X1 OAI21X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_3052_), .B(raddr1_0_bF_buf2_), .C(_3053_), .Y(_3054_) );
MUX2X1 MUX2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_3054_), .B(regs_30__12_), .S(raddr1_1_bF_buf5_), .Y(_3055_) );
NAND2X1 NAND2X1_458 ( .gnd(gnd), .vdd(vdd), .A(regs_26__12_), .B(raddr1_0_bF_buf1_), .Y(_3056_) );
OAI21X1 OAI21X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_1167_), .B(raddr1_0_bF_buf0_), .C(_3056_), .Y(_3057_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(regs_25__12_), .Y(_3058_) );
NAND2X1 NAND2X1_459 ( .gnd(gnd), .vdd(vdd), .A(regs_24__12_), .B(raddr1_0_bF_buf96_), .Y(_3059_) );
OAI21X1 OAI21X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_3058_), .B(raddr1_0_bF_buf95_), .C(_3059_), .Y(_3060_) );
MUX2X1 MUX2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_3060_), .B(_3057_), .S(raddr1_1_bF_buf4_), .Y(_3061_) );
MUX2X1 MUX2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_3061_), .B(_3055_), .S(raddr1_2_bF_buf1_), .Y(_3062_) );
MUX2X1 MUX2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_3062_), .B(_3051_), .S(_2398__bF_buf1), .Y(_3063_) );
MUX2X1 MUX2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_3039_), .B(_3063_), .S(raddr1_4_bF_buf2_), .Y(_5511__12_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(regs_5__13_), .Y(_3064_) );
OAI21X1 OAI21X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_3064_), .B(raddr1_0_bF_buf94_), .C(raddr1_1_bF_buf3_), .Y(_3065_) );
AOI21X1 AOI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(regs_4__13_), .B(raddr1_0_bF_buf93_), .C(_3065_), .Y(_3066_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(regs_6__13_), .B(raddr1_0_bF_buf92_), .Y(_3067_) );
OAI21X1 OAI21X1_1266 ( .gnd(gnd), .vdd(vdd), .A(_2127_), .B(raddr1_0_bF_buf91_), .C(_2415__bF_buf8), .Y(_3068_) );
OAI21X1 OAI21X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_3068_), .B(_3067_), .C(_2399__bF_buf0), .Y(_3069_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(regs_1__13_), .Y(_3070_) );
OAI21X1 OAI21X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_3070_), .B(raddr1_0_bF_buf90_), .C(raddr1_1_bF_buf2_), .Y(_3071_) );
AOI21X1 AOI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(regs_0__13_), .B(raddr1_0_bF_buf89_), .C(_3071_), .Y(_3072_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(regs_3__13_), .Y(_3073_) );
NOR2X1 NOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf88_), .B(_3073_), .Y(_3074_) );
NAND2X1 NAND2X1_460 ( .gnd(gnd), .vdd(vdd), .A(regs_2__13_), .B(raddr1_0_bF_buf87_), .Y(_3075_) );
NAND2X1 NAND2X1_461 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf7), .B(_3075_), .Y(_3076_) );
OAI21X1 OAI21X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_3076_), .B(_3074_), .C(raddr1_2_bF_buf0_), .Y(_3077_) );
OAI22X1 OAI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_3072_), .B(_3077_), .C(_3069_), .D(_3066_), .Y(_3078_) );
NAND2X1 NAND2X1_462 ( .gnd(gnd), .vdd(vdd), .A(regs_10__13_), .B(raddr1_0_bF_buf86_), .Y(_3079_) );
OAI21X1 OAI21X1_1270 ( .gnd(gnd), .vdd(vdd), .A(_1928_), .B(raddr1_0_bF_buf85_), .C(_3079_), .Y(_3080_) );
NAND2X1 NAND2X1_463 ( .gnd(gnd), .vdd(vdd), .A(regs_8__13_), .B(raddr1_0_bF_buf84_), .Y(_3081_) );
OAI21X1 OAI21X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_2026_), .B(raddr1_0_bF_buf83_), .C(_3081_), .Y(_3082_) );
MUX2X1 MUX2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_3082_), .B(_3080_), .S(raddr1_1_bF_buf1_), .Y(_3083_) );
NAND2X1 NAND2X1_464 ( .gnd(gnd), .vdd(vdd), .A(regs_14__13_), .B(raddr1_0_bF_buf82_), .Y(_3084_) );
OAI21X1 OAI21X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_1731_), .B(raddr1_0_bF_buf81_), .C(_3084_), .Y(_3085_) );
NAND2X1 NAND2X1_465 ( .gnd(gnd), .vdd(vdd), .A(regs_12__13_), .B(raddr1_0_bF_buf80_), .Y(_3086_) );
OAI21X1 OAI21X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_1829_), .B(raddr1_0_bF_buf79_), .C(_3086_), .Y(_3087_) );
MUX2X1 MUX2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_3087_), .B(_3085_), .S(raddr1_1_bF_buf0_), .Y(_3088_) );
MUX2X1 MUX2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_3088_), .B(_3083_), .S(_2399__bF_buf8), .Y(_3089_) );
MUX2X1 MUX2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_3089_), .B(_3078_), .S(_2398__bF_buf0), .Y(_3090_) );
OAI21X1 OAI21X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .B(raddr1_0_bF_buf78_), .C(raddr1_1_bF_buf14_bF_buf0_), .Y(_3091_) );
AOI21X1 AOI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(regs_16__13_), .B(raddr1_0_bF_buf77_), .C(_3091_), .Y(_3092_) );
NOR2X1 NOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf76_), .B(_1533_), .Y(_3093_) );
NAND2X1 NAND2X1_466 ( .gnd(gnd), .vdd(vdd), .A(regs_18__13_), .B(raddr1_0_bF_buf75_), .Y(_3094_) );
NAND2X1 NAND2X1_467 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf6), .B(_3094_), .Y(_3095_) );
OAI21X1 OAI21X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_3095_), .B(_3093_), .C(raddr1_2_bF_buf10_), .Y(_3096_) );
OAI21X1 OAI21X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_1434_), .B(raddr1_0_bF_buf74_), .C(raddr1_1_bF_buf13_bF_buf0_), .Y(_3097_) );
AOI21X1 AOI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(regs_20__13_), .B(raddr1_0_bF_buf73_), .C(_3097_), .Y(_3098_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(regs_22__13_), .B(raddr1_0_bF_buf72_), .Y(_3099_) );
OAI21X1 OAI21X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_1336_), .B(raddr1_0_bF_buf71_), .C(_2415__bF_buf5), .Y(_3100_) );
OAI21X1 OAI21X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_3100_), .B(_3099_), .C(_2399__bF_buf7), .Y(_3101_) );
OAI22X1 OAI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_3092_), .B(_3096_), .C(_3101_), .D(_3098_), .Y(_3102_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(regs_29__13_), .Y(_3103_) );
NAND2X1 NAND2X1_468 ( .gnd(gnd), .vdd(vdd), .A(regs_28__13_), .B(raddr1_0_bF_buf70_), .Y(_3104_) );
OAI21X1 OAI21X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_3103_), .B(raddr1_0_bF_buf69_), .C(_3104_), .Y(_3105_) );
MUX2X1 MUX2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_3105_), .B(regs_30__13_), .S(raddr1_1_bF_buf12_bF_buf0_), .Y(_3106_) );
NAND2X1 NAND2X1_469 ( .gnd(gnd), .vdd(vdd), .A(regs_26__13_), .B(raddr1_0_bF_buf68_), .Y(_3107_) );
OAI21X1 OAI21X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(raddr1_0_bF_buf67_), .C(_3107_), .Y(_3108_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(regs_25__13_), .Y(_3109_) );
NAND2X1 NAND2X1_470 ( .gnd(gnd), .vdd(vdd), .A(regs_24__13_), .B(raddr1_0_bF_buf66_), .Y(_3110_) );
OAI21X1 OAI21X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_3109_), .B(raddr1_0_bF_buf65_), .C(_3110_), .Y(_3111_) );
MUX2X1 MUX2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .B(_3108_), .S(raddr1_1_bF_buf11_bF_buf0_), .Y(_3112_) );
MUX2X1 MUX2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_3112_), .B(_3106_), .S(raddr1_2_bF_buf9_), .Y(_3113_) );
MUX2X1 MUX2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_3113_), .B(_3102_), .S(_2398__bF_buf7), .Y(_3114_) );
MUX2X1 MUX2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_3090_), .B(_3114_), .S(raddr1_4_bF_buf1_), .Y(_5511__13_) );
NAND2X1 NAND2X1_471 ( .gnd(gnd), .vdd(vdd), .A(regs_22__14_), .B(raddr1_0_bF_buf64_), .Y(_3115_) );
OAI21X1 OAI21X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_1338_), .B(raddr1_0_bF_buf63_), .C(_3115_), .Y(_3116_) );
NAND2X1 NAND2X1_472 ( .gnd(gnd), .vdd(vdd), .A(regs_20__14_), .B(raddr1_0_bF_buf62_), .Y(_3117_) );
OAI21X1 OAI21X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_1436_), .B(raddr1_0_bF_buf61_), .C(_3117_), .Y(_3118_) );
MUX2X1 MUX2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_3118_), .B(_3116_), .S(raddr1_1_bF_buf10_bF_buf0_), .Y(_3119_) );
NAND2X1 NAND2X1_473 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf6), .B(_3119_), .Y(_3120_) );
NAND2X1 NAND2X1_474 ( .gnd(gnd), .vdd(vdd), .A(regs_18__14_), .B(raddr1_0_bF_buf60_), .Y(_3121_) );
OAI21X1 OAI21X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_1535_), .B(raddr1_0_bF_buf59_), .C(_3121_), .Y(_3122_) );
NAND2X1 NAND2X1_475 ( .gnd(gnd), .vdd(vdd), .A(regs_16__14_), .B(raddr1_0_bF_buf58_), .Y(_3123_) );
OAI21X1 OAI21X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_1633_), .B(raddr1_0_bF_buf57_), .C(_3123_), .Y(_3124_) );
MUX2X1 MUX2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_3124_), .B(_3122_), .S(raddr1_1_bF_buf9_bF_buf0_), .Y(_3125_) );
AOI21X1 AOI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(raddr1_2_bF_buf8_), .B(_3125_), .C(_2398__bF_buf6), .Y(_3126_) );
OAI21X1 OAI21X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_1171_), .B(raddr1_0_bF_buf56_), .C(raddr1_2_bF_buf7_), .Y(_3127_) );
AOI21X1 AOI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(regs_26__14_), .B(raddr1_0_bF_buf55_), .C(_3127_), .Y(_3128_) );
OAI21X1 OAI21X1_1287 ( .gnd(gnd), .vdd(vdd), .A(regs_30__14_), .B(raddr1_2_bF_buf6_), .C(_2415__bF_buf4), .Y(_3129_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(regs_25__14_), .Y(_3130_) );
OAI21X1 OAI21X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_3130_), .B(raddr1_0_bF_buf54_), .C(raddr1_2_bF_buf5_), .Y(_3131_) );
AOI21X1 AOI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(regs_24__14_), .B(raddr1_0_bF_buf53_), .C(_3131_), .Y(_3132_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(regs_29__14_), .Y(_3133_) );
NOR2X1 NOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf52_), .B(_3133_), .Y(_3134_) );
NAND2X1 NAND2X1_476 ( .gnd(gnd), .vdd(vdd), .A(regs_28__14_), .B(raddr1_0_bF_buf51_), .Y(_3135_) );
NAND2X1 NAND2X1_477 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf5), .B(_3135_), .Y(_3136_) );
OAI21X1 OAI21X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_3136_), .B(_3134_), .C(raddr1_1_bF_buf8_), .Y(_3137_) );
OAI22X1 OAI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_3128_), .B(_3129_), .C(_3137_), .D(_3132_), .Y(_3138_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_3138_), .B(_2398__bF_buf5), .C(_3120_), .D(_3126_), .Y(_3139_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(regs_5__14_), .Y(_3140_) );
OAI21X1 OAI21X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_3140_), .B(raddr1_0_bF_buf50_), .C(raddr1_1_bF_buf7_), .Y(_3141_) );
AOI21X1 AOI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(regs_4__14_), .B(raddr1_0_bF_buf49_), .C(_3141_), .Y(_3142_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(regs_6__14_), .B(raddr1_0_bF_buf48_), .Y(_3143_) );
OAI21X1 OAI21X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_2129_), .B(raddr1_0_bF_buf47_), .C(_2415__bF_buf3), .Y(_3144_) );
OAI21X1 OAI21X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_3144_), .B(_3143_), .C(_2399__bF_buf4), .Y(_3145_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(regs_1__14_), .Y(_3146_) );
OAI21X1 OAI21X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_3146_), .B(raddr1_0_bF_buf46_), .C(raddr1_1_bF_buf6_), .Y(_3147_) );
AOI21X1 AOI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(regs_0__14_), .B(raddr1_0_bF_buf45_), .C(_3147_), .Y(_3148_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(regs_3__14_), .Y(_3149_) );
NOR2X1 NOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf44_), .B(_3149_), .Y(_3150_) );
NAND2X1 NAND2X1_478 ( .gnd(gnd), .vdd(vdd), .A(regs_2__14_), .B(raddr1_0_bF_buf43_), .Y(_3151_) );
NAND2X1 NAND2X1_479 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf2), .B(_3151_), .Y(_3152_) );
OAI21X1 OAI21X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_3152_), .B(_3150_), .C(raddr1_2_bF_buf4_), .Y(_3153_) );
OAI22X1 OAI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_3148_), .B(_3153_), .C(_3145_), .D(_3142_), .Y(_3154_) );
NAND2X1 NAND2X1_480 ( .gnd(gnd), .vdd(vdd), .A(regs_10__14_), .B(raddr1_0_bF_buf42_), .Y(_3155_) );
OAI21X1 OAI21X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_1930_), .B(raddr1_0_bF_buf41_), .C(_3155_), .Y(_3156_) );
NAND2X1 NAND2X1_481 ( .gnd(gnd), .vdd(vdd), .A(regs_8__14_), .B(raddr1_0_bF_buf40_), .Y(_3157_) );
OAI21X1 OAI21X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_2028_), .B(raddr1_0_bF_buf39_), .C(_3157_), .Y(_3158_) );
MUX2X1 MUX2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_3158_), .B(_3156_), .S(raddr1_1_bF_buf5_), .Y(_3159_) );
NAND2X1 NAND2X1_482 ( .gnd(gnd), .vdd(vdd), .A(regs_14__14_), .B(raddr1_0_bF_buf38_), .Y(_3160_) );
OAI21X1 OAI21X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_1733_), .B(raddr1_0_bF_buf37_), .C(_3160_), .Y(_3161_) );
NAND2X1 NAND2X1_483 ( .gnd(gnd), .vdd(vdd), .A(regs_12__14_), .B(raddr1_0_bF_buf36_), .Y(_3162_) );
OAI21X1 OAI21X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_1831_), .B(raddr1_0_bF_buf35_), .C(_3162_), .Y(_3163_) );
MUX2X1 MUX2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_3163_), .B(_3161_), .S(raddr1_1_bF_buf4_), .Y(_3164_) );
MUX2X1 MUX2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_3164_), .B(_3159_), .S(_2399__bF_buf3), .Y(_3165_) );
MUX2X1 MUX2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_3165_), .B(_3154_), .S(_2398__bF_buf4), .Y(_3166_) );
MUX2X1 MUX2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_3166_), .B(_3139_), .S(raddr1_4_bF_buf0_), .Y(_5511__14_) );
OAI21X1 OAI21X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_1438_), .B(raddr1_0_bF_buf34_), .C(raddr1_1_bF_buf3_), .Y(_3167_) );
AOI21X1 AOI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(regs_20__15_), .B(raddr1_0_bF_buf33_), .C(_3167_), .Y(_3168_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(regs_22__15_), .B(raddr1_0_bF_buf32_), .Y(_3169_) );
OAI21X1 OAI21X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_1340_), .B(raddr1_0_bF_buf31_), .C(_2415__bF_buf1), .Y(_3170_) );
OAI21X1 OAI21X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_3170_), .B(_3169_), .C(_2399__bF_buf2), .Y(_3171_) );
OAI21X1 OAI21X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .B(raddr1_0_bF_buf30_), .C(raddr1_1_bF_buf2_), .Y(_3172_) );
AOI21X1 AOI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(regs_16__15_), .B(raddr1_0_bF_buf29_), .C(_3172_), .Y(_3173_) );
NOR2X1 NOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf28_), .B(_1537_), .Y(_3174_) );
NAND2X1 NAND2X1_484 ( .gnd(gnd), .vdd(vdd), .A(regs_18__15_), .B(raddr1_0_bF_buf27_), .Y(_3175_) );
NAND2X1 NAND2X1_485 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf0), .B(_3175_), .Y(_3176_) );
OAI21X1 OAI21X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_3176_), .B(_3174_), .C(raddr1_2_bF_buf3_), .Y(_3177_) );
OAI22X1 OAI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_3173_), .B(_3177_), .C(_3171_), .D(_3168_), .Y(_3178_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(regs_29__15_), .Y(_3179_) );
NAND2X1 NAND2X1_486 ( .gnd(gnd), .vdd(vdd), .A(regs_28__15_), .B(raddr1_0_bF_buf26_), .Y(_3180_) );
OAI21X1 OAI21X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_3179_), .B(raddr1_0_bF_buf25_), .C(_3180_), .Y(_3181_) );
MUX2X1 MUX2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_3181_), .B(regs_30__15_), .S(raddr1_1_bF_buf1_), .Y(_3182_) );
NAND2X1 NAND2X1_487 ( .gnd(gnd), .vdd(vdd), .A(regs_26__15_), .B(raddr1_0_bF_buf24_), .Y(_3183_) );
OAI21X1 OAI21X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_1173_), .B(raddr1_0_bF_buf23_), .C(_3183_), .Y(_3184_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(regs_25__15_), .Y(_3185_) );
NAND2X1 NAND2X1_488 ( .gnd(gnd), .vdd(vdd), .A(regs_24__15_), .B(raddr1_0_bF_buf22_), .Y(_3186_) );
OAI21X1 OAI21X1_1306 ( .gnd(gnd), .vdd(vdd), .A(_3185_), .B(raddr1_0_bF_buf21_), .C(_3186_), .Y(_3187_) );
MUX2X1 MUX2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_3187_), .B(_3184_), .S(raddr1_1_bF_buf0_), .Y(_3188_) );
MUX2X1 MUX2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_3188_), .B(_3182_), .S(raddr1_2_bF_buf2_), .Y(_3189_) );
MUX2X1 MUX2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_3189_), .B(_3178_), .S(_2398__bF_buf3), .Y(_3190_) );
NAND2X1 NAND2X1_489 ( .gnd(gnd), .vdd(vdd), .A(regs_6__15_), .B(raddr1_0_bF_buf20_), .Y(_3191_) );
OAI21X1 OAI21X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_2131_), .B(raddr1_0_bF_buf19_), .C(_3191_), .Y(_3192_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(regs_5__15_), .Y(_3193_) );
NAND2X1 NAND2X1_490 ( .gnd(gnd), .vdd(vdd), .A(regs_4__15_), .B(raddr1_0_bF_buf18_), .Y(_3194_) );
OAI21X1 OAI21X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_3193_), .B(raddr1_0_bF_buf17_), .C(_3194_), .Y(_3195_) );
MUX2X1 MUX2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_3195_), .B(_3192_), .S(raddr1_1_bF_buf14_bF_buf3_), .Y(_3196_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(regs_3__15_), .Y(_3197_) );
NAND2X1 NAND2X1_491 ( .gnd(gnd), .vdd(vdd), .A(regs_2__15_), .B(raddr1_0_bF_buf16_), .Y(_3198_) );
OAI21X1 OAI21X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_3197_), .B(raddr1_0_bF_buf15_), .C(_3198_), .Y(_3199_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(regs_1__15_), .Y(_3200_) );
NAND2X1 NAND2X1_492 ( .gnd(gnd), .vdd(vdd), .A(regs_0__15_), .B(raddr1_0_bF_buf14_), .Y(_3201_) );
OAI21X1 OAI21X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_3200_), .B(raddr1_0_bF_buf13_), .C(_3201_), .Y(_3202_) );
MUX2X1 MUX2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_3202_), .B(_3199_), .S(raddr1_1_bF_buf13_bF_buf3_), .Y(_3203_) );
MUX2X1 MUX2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_3203_), .B(_3196_), .S(raddr1_2_bF_buf1_), .Y(_3204_) );
NAND2X1 NAND2X1_493 ( .gnd(gnd), .vdd(vdd), .A(regs_14__15_), .B(raddr1_0_bF_buf12_), .Y(_3205_) );
OAI21X1 OAI21X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .B(raddr1_0_bF_buf11_), .C(_3205_), .Y(_3206_) );
NAND2X1 NAND2X1_494 ( .gnd(gnd), .vdd(vdd), .A(regs_12__15_), .B(raddr1_0_bF_buf10_), .Y(_3207_) );
OAI21X1 OAI21X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_1833_), .B(raddr1_0_bF_buf9_), .C(_3207_), .Y(_3208_) );
MUX2X1 MUX2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_3208_), .B(_3206_), .S(raddr1_1_bF_buf12_bF_buf3_), .Y(_3209_) );
NAND2X1 NAND2X1_495 ( .gnd(gnd), .vdd(vdd), .A(regs_10__15_), .B(raddr1_0_bF_buf8_), .Y(_3210_) );
OAI21X1 OAI21X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_1932_), .B(raddr1_0_bF_buf7_), .C(_3210_), .Y(_3211_) );
NAND2X1 NAND2X1_496 ( .gnd(gnd), .vdd(vdd), .A(regs_8__15_), .B(raddr1_0_bF_buf6_), .Y(_3212_) );
OAI21X1 OAI21X1_1314 ( .gnd(gnd), .vdd(vdd), .A(_2030_), .B(raddr1_0_bF_buf5_), .C(_3212_), .Y(_3213_) );
MUX2X1 MUX2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_3213_), .B(_3211_), .S(raddr1_1_bF_buf11_bF_buf3_), .Y(_3214_) );
MUX2X1 MUX2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_3214_), .B(_3209_), .S(raddr1_2_bF_buf0_), .Y(_3215_) );
MUX2X1 MUX2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_3215_), .B(_3204_), .S(_2398__bF_buf2), .Y(_3216_) );
MUX2X1 MUX2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_3216_), .B(_3190_), .S(raddr1_4_bF_buf4_), .Y(_5511__15_) );
NAND2X1 NAND2X1_497 ( .gnd(gnd), .vdd(vdd), .A(regs_22__16_), .B(raddr1_0_bF_buf4_), .Y(_3217_) );
OAI21X1 OAI21X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_1342_), .B(raddr1_0_bF_buf3_), .C(_3217_), .Y(_3218_) );
NAND2X1 NAND2X1_498 ( .gnd(gnd), .vdd(vdd), .A(regs_20__16_), .B(raddr1_0_bF_buf2_), .Y(_3219_) );
OAI21X1 OAI21X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_1440_), .B(raddr1_0_bF_buf1_), .C(_3219_), .Y(_3220_) );
MUX2X1 MUX2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_3220_), .B(_3218_), .S(raddr1_1_bF_buf10_bF_buf3_), .Y(_3221_) );
NAND2X1 NAND2X1_499 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf1), .B(_3221_), .Y(_3222_) );
NAND2X1 NAND2X1_500 ( .gnd(gnd), .vdd(vdd), .A(regs_18__16_), .B(raddr1_0_bF_buf0_), .Y(_3223_) );
OAI21X1 OAI21X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_1539_), .B(raddr1_0_bF_buf96_), .C(_3223_), .Y(_3224_) );
NAND2X1 NAND2X1_501 ( .gnd(gnd), .vdd(vdd), .A(regs_16__16_), .B(raddr1_0_bF_buf95_), .Y(_3225_) );
OAI21X1 OAI21X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_1637_), .B(raddr1_0_bF_buf94_), .C(_3225_), .Y(_3226_) );
MUX2X1 MUX2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_3224_), .S(raddr1_1_bF_buf9_bF_buf3_), .Y(_3227_) );
AOI21X1 AOI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(raddr1_2_bF_buf10_), .B(_3227_), .C(_2398__bF_buf1), .Y(_3228_) );
OAI21X1 OAI21X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_1175_), .B(raddr1_0_bF_buf93_), .C(raddr1_2_bF_buf9_), .Y(_3229_) );
AOI21X1 AOI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(regs_26__16_), .B(raddr1_0_bF_buf92_), .C(_3229_), .Y(_3230_) );
OAI21X1 OAI21X1_1320 ( .gnd(gnd), .vdd(vdd), .A(regs_30__16_), .B(raddr1_2_bF_buf8_), .C(_2415__bF_buf8), .Y(_3231_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(regs_25__16_), .Y(_3232_) );
OAI21X1 OAI21X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_3232_), .B(raddr1_0_bF_buf91_), .C(raddr1_2_bF_buf7_), .Y(_3233_) );
AOI21X1 AOI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(regs_24__16_), .B(raddr1_0_bF_buf90_), .C(_3233_), .Y(_3234_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(regs_29__16_), .Y(_3235_) );
NOR2X1 NOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf89_), .B(_3235_), .Y(_3236_) );
NAND2X1 NAND2X1_502 ( .gnd(gnd), .vdd(vdd), .A(regs_28__16_), .B(raddr1_0_bF_buf88_), .Y(_3237_) );
NAND2X1 NAND2X1_503 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf0), .B(_3237_), .Y(_3238_) );
OAI21X1 OAI21X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_3238_), .B(_3236_), .C(raddr1_1_bF_buf8_), .Y(_3239_) );
OAI22X1 OAI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_3230_), .B(_3231_), .C(_3239_), .D(_3234_), .Y(_3240_) );
AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_3240_), .B(_2398__bF_buf0), .C(_3222_), .D(_3228_), .Y(_3241_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(regs_5__16_), .Y(_3242_) );
OAI21X1 OAI21X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_3242_), .B(raddr1_0_bF_buf87_), .C(raddr1_1_bF_buf7_), .Y(_3243_) );
AOI21X1 AOI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(regs_4__16_), .B(raddr1_0_bF_buf86_), .C(_3243_), .Y(_3244_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(regs_6__16_), .B(raddr1_0_bF_buf85_), .Y(_3245_) );
OAI21X1 OAI21X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_2133_), .B(raddr1_0_bF_buf84_), .C(_2415__bF_buf7), .Y(_3246_) );
OAI21X1 OAI21X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_3246_), .B(_3245_), .C(_2399__bF_buf8), .Y(_3247_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(regs_1__16_), .Y(_3248_) );
OAI21X1 OAI21X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_3248_), .B(raddr1_0_bF_buf83_), .C(raddr1_1_bF_buf6_), .Y(_3249_) );
AOI21X1 AOI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(regs_0__16_), .B(raddr1_0_bF_buf82_), .C(_3249_), .Y(_3250_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(regs_3__16_), .Y(_3251_) );
NOR2X1 NOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf81_), .B(_3251_), .Y(_3252_) );
NAND2X1 NAND2X1_504 ( .gnd(gnd), .vdd(vdd), .A(regs_2__16_), .B(raddr1_0_bF_buf80_), .Y(_3253_) );
NAND2X1 NAND2X1_505 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf6), .B(_3253_), .Y(_3254_) );
OAI21X1 OAI21X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_3254_), .B(_3252_), .C(raddr1_2_bF_buf6_), .Y(_3255_) );
OAI22X1 OAI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_3250_), .B(_3255_), .C(_3247_), .D(_3244_), .Y(_3256_) );
NAND2X1 NAND2X1_506 ( .gnd(gnd), .vdd(vdd), .A(regs_10__16_), .B(raddr1_0_bF_buf79_), .Y(_3257_) );
OAI21X1 OAI21X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_1934_), .B(raddr1_0_bF_buf78_), .C(_3257_), .Y(_3258_) );
NAND2X1 NAND2X1_507 ( .gnd(gnd), .vdd(vdd), .A(regs_8__16_), .B(raddr1_0_bF_buf77_), .Y(_3259_) );
OAI21X1 OAI21X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_2032_), .B(raddr1_0_bF_buf76_), .C(_3259_), .Y(_3260_) );
MUX2X1 MUX2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_3260_), .B(_3258_), .S(raddr1_1_bF_buf5_), .Y(_3261_) );
NAND2X1 NAND2X1_508 ( .gnd(gnd), .vdd(vdd), .A(regs_14__16_), .B(raddr1_0_bF_buf75_), .Y(_3262_) );
OAI21X1 OAI21X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(raddr1_0_bF_buf74_), .C(_3262_), .Y(_3263_) );
NAND2X1 NAND2X1_509 ( .gnd(gnd), .vdd(vdd), .A(regs_12__16_), .B(raddr1_0_bF_buf73_), .Y(_3264_) );
OAI21X1 OAI21X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_1835_), .B(raddr1_0_bF_buf72_), .C(_3264_), .Y(_3265_) );
MUX2X1 MUX2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_3265_), .B(_3263_), .S(raddr1_1_bF_buf4_), .Y(_3266_) );
MUX2X1 MUX2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_3266_), .B(_3261_), .S(_2399__bF_buf7), .Y(_3267_) );
MUX2X1 MUX2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_3267_), .B(_3256_), .S(_2398__bF_buf7), .Y(_3268_) );
MUX2X1 MUX2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_3268_), .B(_3241_), .S(raddr1_4_bF_buf3_), .Y(_5511__16_) );
NAND2X1 NAND2X1_510 ( .gnd(gnd), .vdd(vdd), .A(regs_22__17_), .B(raddr1_0_bF_buf71_), .Y(_3269_) );
OAI21X1 OAI21X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_1344_), .B(raddr1_0_bF_buf70_), .C(_3269_), .Y(_3270_) );
NAND2X1 NAND2X1_511 ( .gnd(gnd), .vdd(vdd), .A(regs_20__17_), .B(raddr1_0_bF_buf69_), .Y(_3271_) );
OAI21X1 OAI21X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_1442_), .B(raddr1_0_bF_buf68_), .C(_3271_), .Y(_3272_) );
MUX2X1 MUX2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_3272_), .B(_3270_), .S(raddr1_1_bF_buf3_), .Y(_3273_) );
NAND2X1 NAND2X1_512 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf6), .B(_3273_), .Y(_3274_) );
NAND2X1 NAND2X1_513 ( .gnd(gnd), .vdd(vdd), .A(regs_18__17_), .B(raddr1_0_bF_buf67_), .Y(_3275_) );
OAI21X1 OAI21X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_1541_), .B(raddr1_0_bF_buf66_), .C(_3275_), .Y(_3276_) );
NAND2X1 NAND2X1_514 ( .gnd(gnd), .vdd(vdd), .A(regs_16__17_), .B(raddr1_0_bF_buf65_), .Y(_3277_) );
OAI21X1 OAI21X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .B(raddr1_0_bF_buf64_), .C(_3277_), .Y(_3278_) );
MUX2X1 MUX2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_3278_), .B(_3276_), .S(raddr1_1_bF_buf2_), .Y(_3279_) );
AOI21X1 AOI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(raddr1_2_bF_buf5_), .B(_3279_), .C(_2398__bF_buf6), .Y(_3280_) );
OAI21X1 OAI21X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_1177_), .B(raddr1_0_bF_buf63_), .C(raddr1_2_bF_buf4_), .Y(_3281_) );
AOI21X1 AOI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(regs_26__17_), .B(raddr1_0_bF_buf62_), .C(_3281_), .Y(_3282_) );
OAI21X1 OAI21X1_1337 ( .gnd(gnd), .vdd(vdd), .A(regs_30__17_), .B(raddr1_2_bF_buf3_), .C(_2415__bF_buf5), .Y(_3283_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(regs_25__17_), .Y(_3284_) );
OAI21X1 OAI21X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_3284_), .B(raddr1_0_bF_buf61_), .C(raddr1_2_bF_buf2_), .Y(_3285_) );
AOI21X1 AOI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(regs_24__17_), .B(raddr1_0_bF_buf60_), .C(_3285_), .Y(_3286_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(regs_29__17_), .Y(_3287_) );
NOR2X1 NOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf59_), .B(_3287_), .Y(_3288_) );
NAND2X1 NAND2X1_515 ( .gnd(gnd), .vdd(vdd), .A(regs_28__17_), .B(raddr1_0_bF_buf58_), .Y(_3289_) );
NAND2X1 NAND2X1_516 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf5), .B(_3289_), .Y(_3290_) );
OAI21X1 OAI21X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_3290_), .B(_3288_), .C(raddr1_1_bF_buf1_), .Y(_3291_) );
OAI22X1 OAI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(_3282_), .B(_3283_), .C(_3291_), .D(_3286_), .Y(_3292_) );
AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_3292_), .B(_2398__bF_buf5), .C(_3274_), .D(_3280_), .Y(_3293_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(regs_5__17_), .Y(_3294_) );
OAI21X1 OAI21X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_3294_), .B(raddr1_0_bF_buf57_), .C(raddr1_1_bF_buf0_), .Y(_3295_) );
AOI21X1 AOI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(regs_4__17_), .B(raddr1_0_bF_buf56_), .C(_3295_), .Y(_3296_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(regs_6__17_), .B(raddr1_0_bF_buf55_), .Y(_3297_) );
OAI21X1 OAI21X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_2135_), .B(raddr1_0_bF_buf54_), .C(_2415__bF_buf4), .Y(_3298_) );
OAI21X1 OAI21X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_3298_), .B(_3297_), .C(_2399__bF_buf4), .Y(_3299_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(regs_1__17_), .Y(_3300_) );
OAI21X1 OAI21X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_3300_), .B(raddr1_0_bF_buf53_), .C(raddr1_1_bF_buf14_bF_buf2_), .Y(_3301_) );
AOI21X1 AOI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(regs_0__17_), .B(raddr1_0_bF_buf52_), .C(_3301_), .Y(_3302_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(regs_3__17_), .Y(_3303_) );
NOR2X1 NOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf51_), .B(_3303_), .Y(_3304_) );
NAND2X1 NAND2X1_517 ( .gnd(gnd), .vdd(vdd), .A(regs_2__17_), .B(raddr1_0_bF_buf50_), .Y(_3305_) );
NAND2X1 NAND2X1_518 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf3), .B(_3305_), .Y(_3306_) );
OAI21X1 OAI21X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_3306_), .B(_3304_), .C(raddr1_2_bF_buf1_), .Y(_3307_) );
OAI22X1 OAI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_3302_), .B(_3307_), .C(_3299_), .D(_3296_), .Y(_3308_) );
NAND2X1 NAND2X1_519 ( .gnd(gnd), .vdd(vdd), .A(regs_10__17_), .B(raddr1_0_bF_buf49_), .Y(_3309_) );
OAI21X1 OAI21X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_1936_), .B(raddr1_0_bF_buf48_), .C(_3309_), .Y(_3310_) );
NAND2X1 NAND2X1_520 ( .gnd(gnd), .vdd(vdd), .A(regs_8__17_), .B(raddr1_0_bF_buf47_), .Y(_3311_) );
OAI21X1 OAI21X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_2034_), .B(raddr1_0_bF_buf46_), .C(_3311_), .Y(_3312_) );
MUX2X1 MUX2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_3312_), .B(_3310_), .S(raddr1_1_bF_buf13_bF_buf2_), .Y(_3313_) );
NAND2X1 NAND2X1_521 ( .gnd(gnd), .vdd(vdd), .A(regs_14__17_), .B(raddr1_0_bF_buf45_), .Y(_3314_) );
OAI21X1 OAI21X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_1739_), .B(raddr1_0_bF_buf44_), .C(_3314_), .Y(_3315_) );
NAND2X1 NAND2X1_522 ( .gnd(gnd), .vdd(vdd), .A(regs_12__17_), .B(raddr1_0_bF_buf43_), .Y(_3316_) );
OAI21X1 OAI21X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_1837_), .B(raddr1_0_bF_buf42_), .C(_3316_), .Y(_3317_) );
MUX2X1 MUX2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_3317_), .B(_3315_), .S(raddr1_1_bF_buf12_bF_buf2_), .Y(_3318_) );
MUX2X1 MUX2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_3318_), .B(_3313_), .S(_2399__bF_buf3), .Y(_3319_) );
MUX2X1 MUX2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_3319_), .B(_3308_), .S(_2398__bF_buf4), .Y(_3320_) );
MUX2X1 MUX2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_3320_), .B(_3293_), .S(raddr1_4_bF_buf2_), .Y(_5511__17_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(regs_5__18_), .Y(_3321_) );
OAI21X1 OAI21X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_3321_), .B(raddr1_0_bF_buf41_), .C(raddr1_1_bF_buf11_bF_buf2_), .Y(_3322_) );
AOI21X1 AOI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(regs_4__18_), .B(raddr1_0_bF_buf40_), .C(_3322_), .Y(_3323_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(regs_6__18_), .B(raddr1_0_bF_buf39_), .Y(_3324_) );
OAI21X1 OAI21X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_2137_), .B(raddr1_0_bF_buf38_), .C(_2415__bF_buf2), .Y(_3325_) );
OAI21X1 OAI21X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_3325_), .B(_3324_), .C(_2399__bF_buf2), .Y(_3326_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(regs_1__18_), .Y(_3327_) );
OAI21X1 OAI21X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_3327_), .B(raddr1_0_bF_buf37_), .C(raddr1_1_bF_buf10_bF_buf2_), .Y(_3328_) );
AOI21X1 AOI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(regs_0__18_), .B(raddr1_0_bF_buf36_), .C(_3328_), .Y(_3329_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(regs_3__18_), .Y(_3330_) );
NOR2X1 NOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf35_), .B(_3330_), .Y(_3331_) );
NAND2X1 NAND2X1_523 ( .gnd(gnd), .vdd(vdd), .A(regs_2__18_), .B(raddr1_0_bF_buf34_), .Y(_3332_) );
NAND2X1 NAND2X1_524 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf1), .B(_3332_), .Y(_3333_) );
OAI21X1 OAI21X1_1353 ( .gnd(gnd), .vdd(vdd), .A(_3333_), .B(_3331_), .C(raddr1_2_bF_buf0_), .Y(_3334_) );
OAI22X1 OAI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_3329_), .B(_3334_), .C(_3326_), .D(_3323_), .Y(_3335_) );
NAND2X1 NAND2X1_525 ( .gnd(gnd), .vdd(vdd), .A(regs_10__18_), .B(raddr1_0_bF_buf33_), .Y(_3336_) );
OAI21X1 OAI21X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_1938_), .B(raddr1_0_bF_buf32_), .C(_3336_), .Y(_3337_) );
NAND2X1 NAND2X1_526 ( .gnd(gnd), .vdd(vdd), .A(regs_8__18_), .B(raddr1_0_bF_buf31_), .Y(_3338_) );
OAI21X1 OAI21X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_2036_), .B(raddr1_0_bF_buf30_), .C(_3338_), .Y(_3339_) );
MUX2X1 MUX2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_3339_), .B(_3337_), .S(raddr1_1_bF_buf9_bF_buf2_), .Y(_3340_) );
NAND2X1 NAND2X1_527 ( .gnd(gnd), .vdd(vdd), .A(regs_14__18_), .B(raddr1_0_bF_buf29_), .Y(_3341_) );
OAI21X1 OAI21X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_1741_), .B(raddr1_0_bF_buf28_), .C(_3341_), .Y(_3342_) );
NAND2X1 NAND2X1_528 ( .gnd(gnd), .vdd(vdd), .A(regs_12__18_), .B(raddr1_0_bF_buf27_), .Y(_3343_) );
OAI21X1 OAI21X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_1839_), .B(raddr1_0_bF_buf26_), .C(_3343_), .Y(_3344_) );
MUX2X1 MUX2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_3344_), .B(_3342_), .S(raddr1_1_bF_buf8_), .Y(_3345_) );
MUX2X1 MUX2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_3345_), .B(_3340_), .S(_2399__bF_buf1), .Y(_3346_) );
MUX2X1 MUX2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_3346_), .B(_3335_), .S(_2398__bF_buf3), .Y(_3347_) );
OAI21X1 OAI21X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_1641_), .B(raddr1_0_bF_buf25_), .C(raddr1_1_bF_buf7_), .Y(_3348_) );
AOI21X1 AOI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(regs_16__18_), .B(raddr1_0_bF_buf24_), .C(_3348_), .Y(_3349_) );
NOR2X1 NOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf23_), .B(_1543_), .Y(_3350_) );
NAND2X1 NAND2X1_529 ( .gnd(gnd), .vdd(vdd), .A(regs_18__18_), .B(raddr1_0_bF_buf22_), .Y(_3351_) );
NAND2X1 NAND2X1_530 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf0), .B(_3351_), .Y(_3352_) );
OAI21X1 OAI21X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_3352_), .B(_3350_), .C(raddr1_2_bF_buf10_), .Y(_3353_) );
OAI21X1 OAI21X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_1444_), .B(raddr1_0_bF_buf21_), .C(raddr1_1_bF_buf6_), .Y(_3354_) );
AOI21X1 AOI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(regs_20__18_), .B(raddr1_0_bF_buf20_), .C(_3354_), .Y(_3355_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(regs_22__18_), .B(raddr1_0_bF_buf19_), .Y(_3356_) );
OAI21X1 OAI21X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_1346_), .B(raddr1_0_bF_buf18_), .C(_2415__bF_buf8), .Y(_3357_) );
OAI21X1 OAI21X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_3357_), .B(_3356_), .C(_2399__bF_buf0), .Y(_3358_) );
OAI22X1 OAI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_3349_), .B(_3353_), .C(_3358_), .D(_3355_), .Y(_3359_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(regs_29__18_), .Y(_3360_) );
NAND2X1 NAND2X1_531 ( .gnd(gnd), .vdd(vdd), .A(regs_28__18_), .B(raddr1_0_bF_buf17_), .Y(_3361_) );
OAI21X1 OAI21X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_3360_), .B(raddr1_0_bF_buf16_), .C(_3361_), .Y(_3362_) );
MUX2X1 MUX2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_3362_), .B(regs_30__18_), .S(raddr1_1_bF_buf5_), .Y(_3363_) );
NAND2X1 NAND2X1_532 ( .gnd(gnd), .vdd(vdd), .A(regs_26__18_), .B(raddr1_0_bF_buf15_), .Y(_3364_) );
OAI21X1 OAI21X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_1179_), .B(raddr1_0_bF_buf14_), .C(_3364_), .Y(_3365_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(regs_25__18_), .Y(_3366_) );
NAND2X1 NAND2X1_533 ( .gnd(gnd), .vdd(vdd), .A(regs_24__18_), .B(raddr1_0_bF_buf13_), .Y(_3367_) );
OAI21X1 OAI21X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_3366_), .B(raddr1_0_bF_buf12_), .C(_3367_), .Y(_3368_) );
MUX2X1 MUX2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_3368_), .B(_3365_), .S(raddr1_1_bF_buf4_), .Y(_3369_) );
MUX2X1 MUX2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(_3363_), .S(raddr1_2_bF_buf9_), .Y(_3370_) );
MUX2X1 MUX2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_3370_), .B(_3359_), .S(_2398__bF_buf2), .Y(_3371_) );
MUX2X1 MUX2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_3347_), .B(_3371_), .S(raddr1_4_bF_buf1_), .Y(_5511__18_) );
NAND2X1 NAND2X1_534 ( .gnd(gnd), .vdd(vdd), .A(regs_22__19_), .B(raddr1_0_bF_buf11_), .Y(_3372_) );
OAI21X1 OAI21X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_1348_), .B(raddr1_0_bF_buf10_), .C(_3372_), .Y(_3373_) );
NAND2X1 NAND2X1_535 ( .gnd(gnd), .vdd(vdd), .A(regs_20__19_), .B(raddr1_0_bF_buf9_), .Y(_3374_) );
OAI21X1 OAI21X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_1446_), .B(raddr1_0_bF_buf8_), .C(_3374_), .Y(_3375_) );
MUX2X1 MUX2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_3375_), .B(_3373_), .S(raddr1_1_bF_buf3_), .Y(_3376_) );
NAND2X1 NAND2X1_536 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf8), .B(_3376_), .Y(_3377_) );
NAND2X1 NAND2X1_537 ( .gnd(gnd), .vdd(vdd), .A(regs_18__19_), .B(raddr1_0_bF_buf7_), .Y(_3378_) );
OAI21X1 OAI21X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_1545_), .B(raddr1_0_bF_buf6_), .C(_3378_), .Y(_3379_) );
NAND2X1 NAND2X1_538 ( .gnd(gnd), .vdd(vdd), .A(regs_16__19_), .B(raddr1_0_bF_buf5_), .Y(_3380_) );
OAI21X1 OAI21X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .B(raddr1_0_bF_buf4_), .C(_3380_), .Y(_3381_) );
MUX2X1 MUX2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_3381_), .B(_3379_), .S(raddr1_1_bF_buf2_), .Y(_3382_) );
AOI21X1 AOI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(raddr1_2_bF_buf8_), .B(_3382_), .C(_2398__bF_buf1), .Y(_3383_) );
OAI21X1 OAI21X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_1181_), .B(raddr1_0_bF_buf3_), .C(raddr1_2_bF_buf7_), .Y(_3384_) );
AOI21X1 AOI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(regs_26__19_), .B(raddr1_0_bF_buf2_), .C(_3384_), .Y(_3385_) );
OAI21X1 OAI21X1_1371 ( .gnd(gnd), .vdd(vdd), .A(regs_30__19_), .B(raddr1_2_bF_buf6_), .C(_2415__bF_buf7), .Y(_3386_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(regs_25__19_), .Y(_3387_) );
OAI21X1 OAI21X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .B(raddr1_0_bF_buf1_), .C(raddr1_2_bF_buf5_), .Y(_3388_) );
AOI21X1 AOI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(regs_24__19_), .B(raddr1_0_bF_buf0_), .C(_3388_), .Y(_3389_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(regs_29__19_), .Y(_3390_) );
NOR2X1 NOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf96_), .B(_3390_), .Y(_3391_) );
NAND2X1 NAND2X1_539 ( .gnd(gnd), .vdd(vdd), .A(regs_28__19_), .B(raddr1_0_bF_buf95_), .Y(_3392_) );
NAND2X1 NAND2X1_540 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf7), .B(_3392_), .Y(_3393_) );
OAI21X1 OAI21X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_3393_), .B(_3391_), .C(raddr1_1_bF_buf1_), .Y(_3394_) );
OAI22X1 OAI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_3385_), .B(_3386_), .C(_3394_), .D(_3389_), .Y(_3395_) );
AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_3395_), .B(_2398__bF_buf0), .C(_3377_), .D(_3383_), .Y(_3396_) );
NAND2X1 NAND2X1_541 ( .gnd(gnd), .vdd(vdd), .A(regs_6__19_), .B(raddr1_0_bF_buf94_), .Y(_3397_) );
OAI21X1 OAI21X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_2139_), .B(raddr1_0_bF_buf93_), .C(_3397_), .Y(_3398_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(regs_5__19_), .Y(_3399_) );
NAND2X1 NAND2X1_542 ( .gnd(gnd), .vdd(vdd), .A(regs_4__19_), .B(raddr1_0_bF_buf92_), .Y(_3400_) );
OAI21X1 OAI21X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_3399_), .B(raddr1_0_bF_buf91_), .C(_3400_), .Y(_3401_) );
MUX2X1 MUX2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_3401_), .B(_3398_), .S(raddr1_1_bF_buf0_), .Y(_3402_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(regs_3__19_), .Y(_3403_) );
NAND2X1 NAND2X1_543 ( .gnd(gnd), .vdd(vdd), .A(regs_2__19_), .B(raddr1_0_bF_buf90_), .Y(_3404_) );
OAI21X1 OAI21X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_3403_), .B(raddr1_0_bF_buf89_), .C(_3404_), .Y(_3405_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(regs_1__19_), .Y(_3406_) );
NAND2X1 NAND2X1_544 ( .gnd(gnd), .vdd(vdd), .A(regs_0__19_), .B(raddr1_0_bF_buf88_), .Y(_3407_) );
OAI21X1 OAI21X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_3406_), .B(raddr1_0_bF_buf87_), .C(_3407_), .Y(_3408_) );
MUX2X1 MUX2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_3408_), .B(_3405_), .S(raddr1_1_bF_buf14_bF_buf1_), .Y(_3409_) );
MUX2X1 MUX2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_3409_), .B(_3402_), .S(raddr1_2_bF_buf4_), .Y(_3410_) );
NAND2X1 NAND2X1_545 ( .gnd(gnd), .vdd(vdd), .A(regs_10__19_), .B(raddr1_0_bF_buf86_), .Y(_3411_) );
OAI21X1 OAI21X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_1940_), .B(raddr1_0_bF_buf85_), .C(_3411_), .Y(_3412_) );
NAND2X1 NAND2X1_546 ( .gnd(gnd), .vdd(vdd), .A(regs_8__19_), .B(raddr1_0_bF_buf84_), .Y(_3413_) );
OAI21X1 OAI21X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_2038_), .B(raddr1_0_bF_buf83_), .C(_3413_), .Y(_3414_) );
MUX2X1 MUX2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_3414_), .B(_3412_), .S(raddr1_1_bF_buf13_bF_buf1_), .Y(_3415_) );
NAND2X1 NAND2X1_547 ( .gnd(gnd), .vdd(vdd), .A(regs_14__19_), .B(raddr1_0_bF_buf82_), .Y(_3416_) );
OAI21X1 OAI21X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_1743_), .B(raddr1_0_bF_buf81_), .C(_3416_), .Y(_3417_) );
NAND2X1 NAND2X1_548 ( .gnd(gnd), .vdd(vdd), .A(regs_12__19_), .B(raddr1_0_bF_buf80_), .Y(_3418_) );
OAI21X1 OAI21X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_1841_), .B(raddr1_0_bF_buf79_), .C(_3418_), .Y(_3419_) );
MUX2X1 MUX2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_3419_), .B(_3417_), .S(raddr1_1_bF_buf12_bF_buf1_), .Y(_3420_) );
MUX2X1 MUX2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_3420_), .B(_3415_), .S(_2399__bF_buf6), .Y(_3421_) );
MUX2X1 MUX2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_3421_), .B(_3410_), .S(_2398__bF_buf7), .Y(_3422_) );
MUX2X1 MUX2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_3422_), .B(_3396_), .S(raddr1_4_bF_buf0_), .Y(_5511__19_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(regs_5__20_), .Y(_3423_) );
OAI21X1 OAI21X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_3423_), .B(raddr1_0_bF_buf78_), .C(raddr1_1_bF_buf11_bF_buf1_), .Y(_3424_) );
AOI21X1 AOI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(regs_4__20_), .B(raddr1_0_bF_buf77_), .C(_3424_), .Y(_3425_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(regs_6__20_), .B(raddr1_0_bF_buf76_), .Y(_3426_) );
OAI21X1 OAI21X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_2141_), .B(raddr1_0_bF_buf75_), .C(_2415__bF_buf6), .Y(_3427_) );
OAI21X1 OAI21X1_1384 ( .gnd(gnd), .vdd(vdd), .A(_3427_), .B(_3426_), .C(_2399__bF_buf5), .Y(_3428_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(regs_1__20_), .Y(_3429_) );
OAI21X1 OAI21X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_3429_), .B(raddr1_0_bF_buf74_), .C(raddr1_1_bF_buf10_bF_buf1_), .Y(_3430_) );
AOI21X1 AOI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(regs_0__20_), .B(raddr1_0_bF_buf73_), .C(_3430_), .Y(_3431_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(regs_3__20_), .Y(_3432_) );
NOR2X1 NOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf72_), .B(_3432_), .Y(_3433_) );
NAND2X1 NAND2X1_549 ( .gnd(gnd), .vdd(vdd), .A(regs_2__20_), .B(raddr1_0_bF_buf71_), .Y(_3434_) );
NAND2X1 NAND2X1_550 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf5), .B(_3434_), .Y(_3435_) );
OAI21X1 OAI21X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_3435_), .B(_3433_), .C(raddr1_2_bF_buf3_), .Y(_3436_) );
OAI22X1 OAI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_3431_), .B(_3436_), .C(_3428_), .D(_3425_), .Y(_3437_) );
NAND2X1 NAND2X1_551 ( .gnd(gnd), .vdd(vdd), .A(regs_10__20_), .B(raddr1_0_bF_buf70_), .Y(_3438_) );
OAI21X1 OAI21X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_1942_), .B(raddr1_0_bF_buf69_), .C(_3438_), .Y(_3439_) );
NAND2X1 NAND2X1_552 ( .gnd(gnd), .vdd(vdd), .A(regs_8__20_), .B(raddr1_0_bF_buf68_), .Y(_3440_) );
OAI21X1 OAI21X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_2040_), .B(raddr1_0_bF_buf67_), .C(_3440_), .Y(_3441_) );
MUX2X1 MUX2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_3441_), .B(_3439_), .S(raddr1_1_bF_buf9_bF_buf1_), .Y(_3442_) );
NAND2X1 NAND2X1_553 ( .gnd(gnd), .vdd(vdd), .A(regs_14__20_), .B(raddr1_0_bF_buf66_), .Y(_3443_) );
OAI21X1 OAI21X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_1745_), .B(raddr1_0_bF_buf65_), .C(_3443_), .Y(_3444_) );
NAND2X1 NAND2X1_554 ( .gnd(gnd), .vdd(vdd), .A(regs_12__20_), .B(raddr1_0_bF_buf64_), .Y(_3445_) );
OAI21X1 OAI21X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_1843_), .B(raddr1_0_bF_buf63_), .C(_3445_), .Y(_3446_) );
MUX2X1 MUX2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_3446_), .B(_3444_), .S(raddr1_1_bF_buf8_), .Y(_3447_) );
MUX2X1 MUX2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_3447_), .B(_3442_), .S(_2399__bF_buf4), .Y(_3448_) );
MUX2X1 MUX2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_3448_), .B(_3437_), .S(_2398__bF_buf6), .Y(_3449_) );
OAI21X1 OAI21X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_1645_), .B(raddr1_0_bF_buf62_), .C(raddr1_1_bF_buf7_), .Y(_3450_) );
AOI21X1 AOI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(regs_16__20_), .B(raddr1_0_bF_buf61_), .C(_3450_), .Y(_3451_) );
NOR2X1 NOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf60_), .B(_1547_), .Y(_3452_) );
NAND2X1 NAND2X1_555 ( .gnd(gnd), .vdd(vdd), .A(regs_18__20_), .B(raddr1_0_bF_buf59_), .Y(_3453_) );
NAND2X1 NAND2X1_556 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf4), .B(_3453_), .Y(_3454_) );
OAI21X1 OAI21X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_3454_), .B(_3452_), .C(raddr1_2_bF_buf2_), .Y(_3455_) );
OAI21X1 OAI21X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_1448_), .B(raddr1_0_bF_buf58_), .C(raddr1_1_bF_buf6_), .Y(_3456_) );
AOI21X1 AOI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(regs_20__20_), .B(raddr1_0_bF_buf57_), .C(_3456_), .Y(_3457_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(regs_22__20_), .B(raddr1_0_bF_buf56_), .Y(_3458_) );
OAI21X1 OAI21X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_1350_), .B(raddr1_0_bF_buf55_), .C(_2415__bF_buf3), .Y(_3459_) );
OAI21X1 OAI21X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_3459_), .B(_3458_), .C(_2399__bF_buf3), .Y(_3460_) );
OAI22X1 OAI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_3451_), .B(_3455_), .C(_3460_), .D(_3457_), .Y(_3461_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(regs_29__20_), .Y(_3462_) );
NAND2X1 NAND2X1_557 ( .gnd(gnd), .vdd(vdd), .A(regs_28__20_), .B(raddr1_0_bF_buf54_), .Y(_3463_) );
OAI21X1 OAI21X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_3462_), .B(raddr1_0_bF_buf53_), .C(_3463_), .Y(_3464_) );
MUX2X1 MUX2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_3464_), .B(regs_30__20_), .S(raddr1_1_bF_buf5_), .Y(_3465_) );
NAND2X1 NAND2X1_558 ( .gnd(gnd), .vdd(vdd), .A(regs_26__20_), .B(raddr1_0_bF_buf52_), .Y(_3466_) );
OAI21X1 OAI21X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_1183_), .B(raddr1_0_bF_buf51_), .C(_3466_), .Y(_3467_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(regs_25__20_), .Y(_3468_) );
NAND2X1 NAND2X1_559 ( .gnd(gnd), .vdd(vdd), .A(regs_24__20_), .B(raddr1_0_bF_buf50_), .Y(_3469_) );
OAI21X1 OAI21X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_3468_), .B(raddr1_0_bF_buf49_), .C(_3469_), .Y(_3470_) );
MUX2X1 MUX2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_3470_), .B(_3467_), .S(raddr1_1_bF_buf4_), .Y(_3471_) );
MUX2X1 MUX2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_3471_), .B(_3465_), .S(raddr1_2_bF_buf1_), .Y(_3472_) );
MUX2X1 MUX2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_3472_), .B(_3461_), .S(_2398__bF_buf5), .Y(_3473_) );
MUX2X1 MUX2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_3449_), .B(_3473_), .S(raddr1_4_bF_buf4_), .Y(_5511__20_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(regs_5__21_), .Y(_3474_) );
OAI21X1 OAI21X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_3474_), .B(raddr1_0_bF_buf48_), .C(raddr1_1_bF_buf3_), .Y(_3475_) );
AOI21X1 AOI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(regs_4__21_), .B(raddr1_0_bF_buf47_), .C(_3475_), .Y(_3476_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(regs_6__21_), .B(raddr1_0_bF_buf46_), .Y(_3477_) );
OAI21X1 OAI21X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_2143_), .B(raddr1_0_bF_buf45_), .C(_2415__bF_buf2), .Y(_3478_) );
OAI21X1 OAI21X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_3478_), .B(_3477_), .C(_2399__bF_buf2), .Y(_3479_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(regs_1__21_), .Y(_3480_) );
OAI21X1 OAI21X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_3480_), .B(raddr1_0_bF_buf44_), .C(raddr1_1_bF_buf2_), .Y(_3481_) );
AOI21X1 AOI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(regs_0__21_), .B(raddr1_0_bF_buf43_), .C(_3481_), .Y(_3482_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(regs_3__21_), .Y(_3483_) );
NOR2X1 NOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf42_), .B(_3483_), .Y(_3484_) );
NAND2X1 NAND2X1_560 ( .gnd(gnd), .vdd(vdd), .A(regs_2__21_), .B(raddr1_0_bF_buf41_), .Y(_3485_) );
NAND2X1 NAND2X1_561 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf1), .B(_3485_), .Y(_3486_) );
OAI21X1 OAI21X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_3486_), .B(_3484_), .C(raddr1_2_bF_buf0_), .Y(_3487_) );
OAI22X1 OAI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_3482_), .B(_3487_), .C(_3479_), .D(_3476_), .Y(_3488_) );
NAND2X1 NAND2X1_562 ( .gnd(gnd), .vdd(vdd), .A(regs_10__21_), .B(raddr1_0_bF_buf40_), .Y(_3489_) );
OAI21X1 OAI21X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_1944_), .B(raddr1_0_bF_buf39_), .C(_3489_), .Y(_3490_) );
NAND2X1 NAND2X1_563 ( .gnd(gnd), .vdd(vdd), .A(regs_8__21_), .B(raddr1_0_bF_buf38_), .Y(_3491_) );
OAI21X1 OAI21X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_2042_), .B(raddr1_0_bF_buf37_), .C(_3491_), .Y(_3492_) );
MUX2X1 MUX2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_3492_), .B(_3490_), .S(raddr1_1_bF_buf1_), .Y(_3493_) );
NAND2X1 NAND2X1_564 ( .gnd(gnd), .vdd(vdd), .A(regs_14__21_), .B(raddr1_0_bF_buf36_), .Y(_3494_) );
OAI21X1 OAI21X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_1747_), .B(raddr1_0_bF_buf35_), .C(_3494_), .Y(_3495_) );
NAND2X1 NAND2X1_565 ( .gnd(gnd), .vdd(vdd), .A(regs_12__21_), .B(raddr1_0_bF_buf34_), .Y(_3496_) );
OAI21X1 OAI21X1_1407 ( .gnd(gnd), .vdd(vdd), .A(_1845_), .B(raddr1_0_bF_buf33_), .C(_3496_), .Y(_3497_) );
MUX2X1 MUX2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_3497_), .B(_3495_), .S(raddr1_1_bF_buf0_), .Y(_3498_) );
MUX2X1 MUX2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_3498_), .B(_3493_), .S(_2399__bF_buf1), .Y(_3499_) );
MUX2X1 MUX2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_3499_), .B(_3488_), .S(_2398__bF_buf4), .Y(_3500_) );
OAI21X1 OAI21X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_1647_), .B(raddr1_0_bF_buf32_), .C(raddr1_1_bF_buf14_bF_buf0_), .Y(_3501_) );
AOI21X1 AOI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(regs_16__21_), .B(raddr1_0_bF_buf31_), .C(_3501_), .Y(_3502_) );
NOR2X1 NOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf30_), .B(_1549_), .Y(_3503_) );
NAND2X1 NAND2X1_566 ( .gnd(gnd), .vdd(vdd), .A(regs_18__21_), .B(raddr1_0_bF_buf29_), .Y(_3504_) );
NAND2X1 NAND2X1_567 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf0), .B(_3504_), .Y(_3505_) );
OAI21X1 OAI21X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_3505_), .B(_3503_), .C(raddr1_2_bF_buf10_), .Y(_3506_) );
OAI21X1 OAI21X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_1450_), .B(raddr1_0_bF_buf28_), .C(raddr1_1_bF_buf13_bF_buf0_), .Y(_3507_) );
AOI21X1 AOI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(regs_20__21_), .B(raddr1_0_bF_buf27_), .C(_3507_), .Y(_3508_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(regs_22__21_), .B(raddr1_0_bF_buf26_), .Y(_3509_) );
OAI21X1 OAI21X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_1352_), .B(raddr1_0_bF_buf25_), .C(_2415__bF_buf8), .Y(_3510_) );
OAI21X1 OAI21X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_3510_), .B(_3509_), .C(_2399__bF_buf0), .Y(_3511_) );
OAI22X1 OAI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_3502_), .B(_3506_), .C(_3511_), .D(_3508_), .Y(_3512_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(regs_29__21_), .Y(_3513_) );
NAND2X1 NAND2X1_568 ( .gnd(gnd), .vdd(vdd), .A(regs_28__21_), .B(raddr1_0_bF_buf24_), .Y(_3514_) );
OAI21X1 OAI21X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_3513_), .B(raddr1_0_bF_buf23_), .C(_3514_), .Y(_3515_) );
MUX2X1 MUX2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_3515_), .B(regs_30__21_), .S(raddr1_1_bF_buf12_bF_buf0_), .Y(_3516_) );
NAND2X1 NAND2X1_569 ( .gnd(gnd), .vdd(vdd), .A(regs_26__21_), .B(raddr1_0_bF_buf22_), .Y(_3517_) );
OAI21X1 OAI21X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_1185_), .B(raddr1_0_bF_buf21_), .C(_3517_), .Y(_3518_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(regs_25__21_), .Y(_3519_) );
NAND2X1 NAND2X1_570 ( .gnd(gnd), .vdd(vdd), .A(regs_24__21_), .B(raddr1_0_bF_buf20_), .Y(_3520_) );
OAI21X1 OAI21X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_3519_), .B(raddr1_0_bF_buf19_), .C(_3520_), .Y(_3521_) );
MUX2X1 MUX2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_3521_), .B(_3518_), .S(raddr1_1_bF_buf11_bF_buf0_), .Y(_3522_) );
MUX2X1 MUX2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_3522_), .B(_3516_), .S(raddr1_2_bF_buf9_), .Y(_3523_) );
MUX2X1 MUX2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_3523_), .B(_3512_), .S(_2398__bF_buf3), .Y(_3524_) );
MUX2X1 MUX2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_3500_), .B(_3524_), .S(raddr1_4_bF_buf3_), .Y(_5511__21_) );
OAI21X1 OAI21X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_1452_), .B(raddr1_0_bF_buf18_), .C(raddr1_1_bF_buf10_bF_buf0_), .Y(_3525_) );
AOI21X1 AOI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(regs_20__22_), .B(raddr1_0_bF_buf17_), .C(_3525_), .Y(_3526_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(regs_22__22_), .B(raddr1_0_bF_buf16_), .Y(_3527_) );
OAI21X1 OAI21X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_1354_), .B(raddr1_0_bF_buf15_), .C(_2415__bF_buf7), .Y(_3528_) );
OAI21X1 OAI21X1_1418 ( .gnd(gnd), .vdd(vdd), .A(_3528_), .B(_3527_), .C(_2399__bF_buf8), .Y(_3529_) );
OAI21X1 OAI21X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_1649_), .B(raddr1_0_bF_buf14_), .C(raddr1_1_bF_buf9_bF_buf0_), .Y(_3530_) );
AOI21X1 AOI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(regs_16__22_), .B(raddr1_0_bF_buf13_), .C(_3530_), .Y(_3531_) );
NOR2X1 NOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf12_), .B(_1551_), .Y(_3532_) );
NAND2X1 NAND2X1_571 ( .gnd(gnd), .vdd(vdd), .A(regs_18__22_), .B(raddr1_0_bF_buf11_), .Y(_3533_) );
NAND2X1 NAND2X1_572 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf6), .B(_3533_), .Y(_3534_) );
OAI21X1 OAI21X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_3534_), .B(_3532_), .C(raddr1_2_bF_buf8_), .Y(_3535_) );
OAI22X1 OAI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_3531_), .B(_3535_), .C(_3529_), .D(_3526_), .Y(_3536_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(regs_29__22_), .Y(_3537_) );
NAND2X1 NAND2X1_573 ( .gnd(gnd), .vdd(vdd), .A(regs_28__22_), .B(raddr1_0_bF_buf10_), .Y(_3538_) );
OAI21X1 OAI21X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_3537_), .B(raddr1_0_bF_buf9_), .C(_3538_), .Y(_3539_) );
MUX2X1 MUX2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_3539_), .B(regs_30__22_), .S(raddr1_1_bF_buf8_), .Y(_3540_) );
NAND2X1 NAND2X1_574 ( .gnd(gnd), .vdd(vdd), .A(regs_26__22_), .B(raddr1_0_bF_buf8_), .Y(_3541_) );
OAI21X1 OAI21X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_1187_), .B(raddr1_0_bF_buf7_), .C(_3541_), .Y(_3542_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(regs_25__22_), .Y(_3543_) );
NAND2X1 NAND2X1_575 ( .gnd(gnd), .vdd(vdd), .A(regs_24__22_), .B(raddr1_0_bF_buf6_), .Y(_3544_) );
OAI21X1 OAI21X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_3543_), .B(raddr1_0_bF_buf5_), .C(_3544_), .Y(_3545_) );
MUX2X1 MUX2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_3545_), .B(_3542_), .S(raddr1_1_bF_buf7_), .Y(_3546_) );
MUX2X1 MUX2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_3546_), .B(_3540_), .S(raddr1_2_bF_buf7_), .Y(_3547_) );
MUX2X1 MUX2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_3547_), .B(_3536_), .S(_2398__bF_buf2), .Y(_3548_) );
NAND2X1 NAND2X1_576 ( .gnd(gnd), .vdd(vdd), .A(regs_6__22_), .B(raddr1_0_bF_buf4_), .Y(_3549_) );
OAI21X1 OAI21X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_2145_), .B(raddr1_0_bF_buf3_), .C(_3549_), .Y(_3550_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(regs_5__22_), .Y(_3551_) );
NAND2X1 NAND2X1_577 ( .gnd(gnd), .vdd(vdd), .A(regs_4__22_), .B(raddr1_0_bF_buf2_), .Y(_3552_) );
OAI21X1 OAI21X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_3551_), .B(raddr1_0_bF_buf1_), .C(_3552_), .Y(_3553_) );
MUX2X1 MUX2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_3553_), .B(_3550_), .S(raddr1_1_bF_buf6_), .Y(_3554_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(regs_3__22_), .Y(_3555_) );
NAND2X1 NAND2X1_578 ( .gnd(gnd), .vdd(vdd), .A(regs_2__22_), .B(raddr1_0_bF_buf0_), .Y(_3556_) );
OAI21X1 OAI21X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_3555_), .B(raddr1_0_bF_buf96_), .C(_3556_), .Y(_3557_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(regs_1__22_), .Y(_3558_) );
NAND2X1 NAND2X1_579 ( .gnd(gnd), .vdd(vdd), .A(regs_0__22_), .B(raddr1_0_bF_buf95_), .Y(_3559_) );
OAI21X1 OAI21X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_3558_), .B(raddr1_0_bF_buf94_), .C(_3559_), .Y(_3560_) );
MUX2X1 MUX2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_3560_), .B(_3557_), .S(raddr1_1_bF_buf5_), .Y(_3561_) );
MUX2X1 MUX2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_3561_), .B(_3554_), .S(raddr1_2_bF_buf6_), .Y(_3562_) );
NAND2X1 NAND2X1_580 ( .gnd(gnd), .vdd(vdd), .A(regs_14__22_), .B(raddr1_0_bF_buf93_), .Y(_3563_) );
OAI21X1 OAI21X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_1749_), .B(raddr1_0_bF_buf92_), .C(_3563_), .Y(_3564_) );
NAND2X1 NAND2X1_581 ( .gnd(gnd), .vdd(vdd), .A(regs_12__22_), .B(raddr1_0_bF_buf91_), .Y(_3565_) );
OAI21X1 OAI21X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_1847_), .B(raddr1_0_bF_buf90_), .C(_3565_), .Y(_3566_) );
MUX2X1 MUX2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_3566_), .B(_3564_), .S(raddr1_1_bF_buf4_), .Y(_3567_) );
NAND2X1 NAND2X1_582 ( .gnd(gnd), .vdd(vdd), .A(regs_10__22_), .B(raddr1_0_bF_buf89_), .Y(_3568_) );
OAI21X1 OAI21X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(raddr1_0_bF_buf88_), .C(_3568_), .Y(_3569_) );
NAND2X1 NAND2X1_583 ( .gnd(gnd), .vdd(vdd), .A(regs_8__22_), .B(raddr1_0_bF_buf87_), .Y(_3570_) );
OAI21X1 OAI21X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_2044_), .B(raddr1_0_bF_buf86_), .C(_3570_), .Y(_3571_) );
MUX2X1 MUX2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_3571_), .B(_3569_), .S(raddr1_1_bF_buf3_), .Y(_3572_) );
MUX2X1 MUX2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_3572_), .B(_3567_), .S(raddr1_2_bF_buf5_), .Y(_3573_) );
MUX2X1 MUX2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_3573_), .B(_3562_), .S(_2398__bF_buf1), .Y(_3574_) );
MUX2X1 MUX2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_3574_), .B(_3548_), .S(raddr1_4_bF_buf2_), .Y(_5511__22_) );
OAI21X1 OAI21X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_1454_), .B(raddr1_0_bF_buf85_), .C(raddr1_1_bF_buf2_), .Y(_3575_) );
AOI21X1 AOI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(regs_20__23_), .B(raddr1_0_bF_buf84_), .C(_3575_), .Y(_3576_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(regs_22__23_), .B(raddr1_0_bF_buf83_), .Y(_3577_) );
OAI21X1 OAI21X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_1356_), .B(raddr1_0_bF_buf82_), .C(_2415__bF_buf5), .Y(_3578_) );
OAI21X1 OAI21X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_3578_), .B(_3577_), .C(_2399__bF_buf7), .Y(_3579_) );
OAI21X1 OAI21X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_1651_), .B(raddr1_0_bF_buf81_), .C(raddr1_1_bF_buf1_), .Y(_3580_) );
AOI21X1 AOI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(regs_16__23_), .B(raddr1_0_bF_buf80_), .C(_3580_), .Y(_3581_) );
NOR2X1 NOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf79_), .B(_1553_), .Y(_3582_) );
NAND2X1 NAND2X1_584 ( .gnd(gnd), .vdd(vdd), .A(regs_18__23_), .B(raddr1_0_bF_buf78_), .Y(_3583_) );
NAND2X1 NAND2X1_585 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf4), .B(_3583_), .Y(_3584_) );
OAI21X1 OAI21X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_3584_), .B(_3582_), .C(raddr1_2_bF_buf4_), .Y(_3585_) );
OAI22X1 OAI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_3581_), .B(_3585_), .C(_3579_), .D(_3576_), .Y(_3586_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(regs_29__23_), .Y(_3587_) );
NAND2X1 NAND2X1_586 ( .gnd(gnd), .vdd(vdd), .A(regs_28__23_), .B(raddr1_0_bF_buf77_), .Y(_3588_) );
OAI21X1 OAI21X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_3587_), .B(raddr1_0_bF_buf76_), .C(_3588_), .Y(_3589_) );
MUX2X1 MUX2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_3589_), .B(regs_30__23_), .S(raddr1_1_bF_buf0_), .Y(_3590_) );
NAND2X1 NAND2X1_587 ( .gnd(gnd), .vdd(vdd), .A(regs_26__23_), .B(raddr1_0_bF_buf75_), .Y(_3591_) );
OAI21X1 OAI21X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_1189_), .B(raddr1_0_bF_buf74_), .C(_3591_), .Y(_3592_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(regs_25__23_), .Y(_3593_) );
NAND2X1 NAND2X1_588 ( .gnd(gnd), .vdd(vdd), .A(regs_24__23_), .B(raddr1_0_bF_buf73_), .Y(_3594_) );
OAI21X1 OAI21X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_3593_), .B(raddr1_0_bF_buf72_), .C(_3594_), .Y(_3595_) );
MUX2X1 MUX2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_3595_), .B(_3592_), .S(raddr1_1_bF_buf14_bF_buf3_), .Y(_3596_) );
MUX2X1 MUX2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_3596_), .B(_3590_), .S(raddr1_2_bF_buf3_), .Y(_3597_) );
MUX2X1 MUX2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_3597_), .B(_3586_), .S(_2398__bF_buf0), .Y(_3598_) );
NAND2X1 NAND2X1_589 ( .gnd(gnd), .vdd(vdd), .A(regs_6__23_), .B(raddr1_0_bF_buf71_), .Y(_3599_) );
OAI21X1 OAI21X1_1440 ( .gnd(gnd), .vdd(vdd), .A(_2147_), .B(raddr1_0_bF_buf70_), .C(_3599_), .Y(_3600_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(regs_5__23_), .Y(_3601_) );
NAND2X1 NAND2X1_590 ( .gnd(gnd), .vdd(vdd), .A(regs_4__23_), .B(raddr1_0_bF_buf69_), .Y(_3602_) );
OAI21X1 OAI21X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_3601_), .B(raddr1_0_bF_buf68_), .C(_3602_), .Y(_3603_) );
MUX2X1 MUX2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_3603_), .B(_3600_), .S(raddr1_1_bF_buf13_bF_buf3_), .Y(_3604_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(regs_3__23_), .Y(_3605_) );
NAND2X1 NAND2X1_591 ( .gnd(gnd), .vdd(vdd), .A(regs_2__23_), .B(raddr1_0_bF_buf67_), .Y(_3606_) );
OAI21X1 OAI21X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_3605_), .B(raddr1_0_bF_buf66_), .C(_3606_), .Y(_3607_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(regs_1__23_), .Y(_3608_) );
NAND2X1 NAND2X1_592 ( .gnd(gnd), .vdd(vdd), .A(regs_0__23_), .B(raddr1_0_bF_buf65_), .Y(_3609_) );
OAI21X1 OAI21X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_3608_), .B(raddr1_0_bF_buf64_), .C(_3609_), .Y(_3610_) );
MUX2X1 MUX2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_3610_), .B(_3607_), .S(raddr1_1_bF_buf12_bF_buf3_), .Y(_3611_) );
MUX2X1 MUX2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_3611_), .B(_3604_), .S(raddr1_2_bF_buf2_), .Y(_3612_) );
NAND2X1 NAND2X1_593 ( .gnd(gnd), .vdd(vdd), .A(regs_14__23_), .B(raddr1_0_bF_buf63_), .Y(_3613_) );
OAI21X1 OAI21X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_1751_), .B(raddr1_0_bF_buf62_), .C(_3613_), .Y(_3614_) );
NAND2X1 NAND2X1_594 ( .gnd(gnd), .vdd(vdd), .A(regs_12__23_), .B(raddr1_0_bF_buf61_), .Y(_3615_) );
OAI21X1 OAI21X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_1849_), .B(raddr1_0_bF_buf60_), .C(_3615_), .Y(_3616_) );
MUX2X1 MUX2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_3616_), .B(_3614_), .S(raddr1_1_bF_buf11_bF_buf3_), .Y(_3617_) );
NAND2X1 NAND2X1_595 ( .gnd(gnd), .vdd(vdd), .A(regs_10__23_), .B(raddr1_0_bF_buf59_), .Y(_3618_) );
OAI21X1 OAI21X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_1948_), .B(raddr1_0_bF_buf58_), .C(_3618_), .Y(_3619_) );
NAND2X1 NAND2X1_596 ( .gnd(gnd), .vdd(vdd), .A(regs_8__23_), .B(raddr1_0_bF_buf57_), .Y(_3620_) );
OAI21X1 OAI21X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_2046_), .B(raddr1_0_bF_buf56_), .C(_3620_), .Y(_3621_) );
MUX2X1 MUX2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_3621_), .B(_3619_), .S(raddr1_1_bF_buf10_bF_buf3_), .Y(_3622_) );
MUX2X1 MUX2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_3622_), .B(_3617_), .S(raddr1_2_bF_buf1_), .Y(_3623_) );
MUX2X1 MUX2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_3623_), .B(_3612_), .S(_2398__bF_buf7), .Y(_3624_) );
MUX2X1 MUX2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_3624_), .B(_3598_), .S(raddr1_4_bF_buf1_), .Y(_5511__23_) );
OAI21X1 OAI21X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_1456_), .B(raddr1_0_bF_buf55_), .C(raddr1_1_bF_buf9_bF_buf3_), .Y(_3625_) );
AOI21X1 AOI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(regs_20__24_), .B(raddr1_0_bF_buf54_), .C(_3625_), .Y(_3626_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(regs_22__24_), .B(raddr1_0_bF_buf53_), .Y(_3627_) );
OAI21X1 OAI21X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_1358_), .B(raddr1_0_bF_buf52_), .C(_2415__bF_buf3), .Y(_3628_) );
OAI21X1 OAI21X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_3628_), .B(_3627_), .C(_2399__bF_buf6), .Y(_3629_) );
OAI21X1 OAI21X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .B(raddr1_0_bF_buf51_), .C(raddr1_1_bF_buf8_), .Y(_3630_) );
AOI21X1 AOI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(regs_16__24_), .B(raddr1_0_bF_buf50_), .C(_3630_), .Y(_3631_) );
NOR2X1 NOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf49_), .B(_1555_), .Y(_3632_) );
NAND2X1 NAND2X1_597 ( .gnd(gnd), .vdd(vdd), .A(regs_18__24_), .B(raddr1_0_bF_buf48_), .Y(_3633_) );
NAND2X1 NAND2X1_598 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf2), .B(_3633_), .Y(_3634_) );
OAI21X1 OAI21X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_3634_), .B(_3632_), .C(raddr1_2_bF_buf0_), .Y(_3635_) );
OAI22X1 OAI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_3631_), .B(_3635_), .C(_3629_), .D(_3626_), .Y(_3636_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(regs_29__24_), .Y(_3637_) );
NAND2X1 NAND2X1_599 ( .gnd(gnd), .vdd(vdd), .A(regs_28__24_), .B(raddr1_0_bF_buf47_), .Y(_3638_) );
OAI21X1 OAI21X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_3637_), .B(raddr1_0_bF_buf46_), .C(_3638_), .Y(_3639_) );
MUX2X1 MUX2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_3639_), .B(regs_30__24_), .S(raddr1_1_bF_buf7_), .Y(_3640_) );
NAND2X1 NAND2X1_600 ( .gnd(gnd), .vdd(vdd), .A(regs_26__24_), .B(raddr1_0_bF_buf45_), .Y(_3641_) );
OAI21X1 OAI21X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_1191_), .B(raddr1_0_bF_buf44_), .C(_3641_), .Y(_3642_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(regs_25__24_), .Y(_3643_) );
NAND2X1 NAND2X1_601 ( .gnd(gnd), .vdd(vdd), .A(regs_24__24_), .B(raddr1_0_bF_buf43_), .Y(_3644_) );
OAI21X1 OAI21X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_3643_), .B(raddr1_0_bF_buf42_), .C(_3644_), .Y(_3645_) );
MUX2X1 MUX2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_3645_), .B(_3642_), .S(raddr1_1_bF_buf6_), .Y(_3646_) );
MUX2X1 MUX2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_3646_), .B(_3640_), .S(raddr1_2_bF_buf10_), .Y(_3647_) );
MUX2X1 MUX2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_3647_), .B(_3636_), .S(_2398__bF_buf6), .Y(_3648_) );
NAND2X1 NAND2X1_602 ( .gnd(gnd), .vdd(vdd), .A(regs_6__24_), .B(raddr1_0_bF_buf41_), .Y(_3649_) );
OAI21X1 OAI21X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_2149_), .B(raddr1_0_bF_buf40_), .C(_3649_), .Y(_3650_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(regs_5__24_), .Y(_3651_) );
NAND2X1 NAND2X1_603 ( .gnd(gnd), .vdd(vdd), .A(regs_4__24_), .B(raddr1_0_bF_buf39_), .Y(_3652_) );
OAI21X1 OAI21X1_1457 ( .gnd(gnd), .vdd(vdd), .A(_3651_), .B(raddr1_0_bF_buf38_), .C(_3652_), .Y(_3653_) );
MUX2X1 MUX2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_3653_), .B(_3650_), .S(raddr1_1_bF_buf5_), .Y(_3654_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(regs_3__24_), .Y(_3655_) );
NAND2X1 NAND2X1_604 ( .gnd(gnd), .vdd(vdd), .A(regs_2__24_), .B(raddr1_0_bF_buf37_), .Y(_3656_) );
OAI21X1 OAI21X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_3655_), .B(raddr1_0_bF_buf36_), .C(_3656_), .Y(_3657_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(regs_1__24_), .Y(_3658_) );
NAND2X1 NAND2X1_605 ( .gnd(gnd), .vdd(vdd), .A(regs_0__24_), .B(raddr1_0_bF_buf35_), .Y(_3659_) );
OAI21X1 OAI21X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_3658_), .B(raddr1_0_bF_buf34_), .C(_3659_), .Y(_3660_) );
MUX2X1 MUX2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_3660_), .B(_3657_), .S(raddr1_1_bF_buf4_), .Y(_3661_) );
MUX2X1 MUX2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_3661_), .B(_3654_), .S(raddr1_2_bF_buf9_), .Y(_3662_) );
NAND2X1 NAND2X1_606 ( .gnd(gnd), .vdd(vdd), .A(regs_10__24_), .B(raddr1_0_bF_buf33_), .Y(_3663_) );
OAI21X1 OAI21X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_1950_), .B(raddr1_0_bF_buf32_), .C(_3663_), .Y(_3664_) );
NAND2X1 NAND2X1_607 ( .gnd(gnd), .vdd(vdd), .A(regs_8__24_), .B(raddr1_0_bF_buf31_), .Y(_3665_) );
OAI21X1 OAI21X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_2048_), .B(raddr1_0_bF_buf30_), .C(_3665_), .Y(_3666_) );
MUX2X1 MUX2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_3666_), .B(_3664_), .S(raddr1_1_bF_buf3_), .Y(_3667_) );
NAND2X1 NAND2X1_608 ( .gnd(gnd), .vdd(vdd), .A(regs_14__24_), .B(raddr1_0_bF_buf29_), .Y(_3668_) );
OAI21X1 OAI21X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_1753_), .B(raddr1_0_bF_buf28_), .C(_3668_), .Y(_3669_) );
NAND2X1 NAND2X1_609 ( .gnd(gnd), .vdd(vdd), .A(regs_12__24_), .B(raddr1_0_bF_buf27_), .Y(_3670_) );
OAI21X1 OAI21X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_1851_), .B(raddr1_0_bF_buf26_), .C(_3670_), .Y(_3671_) );
MUX2X1 MUX2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_3671_), .B(_3669_), .S(raddr1_1_bF_buf2_), .Y(_3672_) );
MUX2X1 MUX2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_3672_), .B(_3667_), .S(_2399__bF_buf5), .Y(_3673_) );
MUX2X1 MUX2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_3673_), .B(_3662_), .S(_2398__bF_buf5), .Y(_3674_) );
MUX2X1 MUX2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_3674_), .B(_3648_), .S(raddr1_4_bF_buf0_), .Y(_5511__24_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(regs_5__25_), .Y(_3675_) );
OAI21X1 OAI21X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_3675_), .B(raddr1_0_bF_buf25_), .C(raddr1_1_bF_buf1_), .Y(_3676_) );
AOI21X1 AOI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(regs_4__25_), .B(raddr1_0_bF_buf24_), .C(_3676_), .Y(_3677_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(regs_6__25_), .B(raddr1_0_bF_buf23_), .Y(_3678_) );
OAI21X1 OAI21X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_2151_), .B(raddr1_0_bF_buf22_), .C(_2415__bF_buf1), .Y(_3679_) );
OAI21X1 OAI21X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_3679_), .B(_3678_), .C(_2399__bF_buf4), .Y(_3680_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(regs_1__25_), .Y(_3681_) );
OAI21X1 OAI21X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_3681_), .B(raddr1_0_bF_buf21_), .C(raddr1_1_bF_buf0_), .Y(_3682_) );
AOI21X1 AOI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(regs_0__25_), .B(raddr1_0_bF_buf20_), .C(_3682_), .Y(_3683_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(regs_3__25_), .Y(_3684_) );
NOR2X1 NOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf19_), .B(_3684_), .Y(_3685_) );
NAND2X1 NAND2X1_610 ( .gnd(gnd), .vdd(vdd), .A(regs_2__25_), .B(raddr1_0_bF_buf18_), .Y(_3686_) );
NAND2X1 NAND2X1_611 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf0), .B(_3686_), .Y(_3687_) );
OAI21X1 OAI21X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_3687_), .B(_3685_), .C(raddr1_2_bF_buf8_), .Y(_3688_) );
OAI22X1 OAI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_3683_), .B(_3688_), .C(_3680_), .D(_3677_), .Y(_3689_) );
NAND2X1 NAND2X1_612 ( .gnd(gnd), .vdd(vdd), .A(regs_10__25_), .B(raddr1_0_bF_buf17_), .Y(_3690_) );
OAI21X1 OAI21X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_1952_), .B(raddr1_0_bF_buf16_), .C(_3690_), .Y(_3691_) );
NAND2X1 NAND2X1_613 ( .gnd(gnd), .vdd(vdd), .A(regs_8__25_), .B(raddr1_0_bF_buf15_), .Y(_3692_) );
OAI21X1 OAI21X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_2050_), .B(raddr1_0_bF_buf14_), .C(_3692_), .Y(_3693_) );
MUX2X1 MUX2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_3693_), .B(_3691_), .S(raddr1_1_bF_buf14_bF_buf2_), .Y(_3694_) );
NAND2X1 NAND2X1_614 ( .gnd(gnd), .vdd(vdd), .A(regs_14__25_), .B(raddr1_0_bF_buf13_), .Y(_3695_) );
OAI21X1 OAI21X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_1755_), .B(raddr1_0_bF_buf12_), .C(_3695_), .Y(_3696_) );
NAND2X1 NAND2X1_615 ( .gnd(gnd), .vdd(vdd), .A(regs_12__25_), .B(raddr1_0_bF_buf11_), .Y(_3697_) );
OAI21X1 OAI21X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_1853_), .B(raddr1_0_bF_buf10_), .C(_3697_), .Y(_3698_) );
MUX2X1 MUX2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_3698_), .B(_3696_), .S(raddr1_1_bF_buf13_bF_buf2_), .Y(_3699_) );
MUX2X1 MUX2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_3699_), .B(_3694_), .S(_2399__bF_buf3), .Y(_3700_) );
MUX2X1 MUX2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_3700_), .B(_3689_), .S(_2398__bF_buf4), .Y(_3701_) );
OAI21X1 OAI21X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .B(raddr1_0_bF_buf9_), .C(raddr1_1_bF_buf12_bF_buf2_), .Y(_3702_) );
AOI21X1 AOI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(regs_16__25_), .B(raddr1_0_bF_buf8_), .C(_3702_), .Y(_3703_) );
NOR2X1 NOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf7_), .B(_1557_), .Y(_3704_) );
NAND2X1 NAND2X1_616 ( .gnd(gnd), .vdd(vdd), .A(regs_18__25_), .B(raddr1_0_bF_buf6_), .Y(_3705_) );
NAND2X1 NAND2X1_617 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf8), .B(_3705_), .Y(_3706_) );
OAI21X1 OAI21X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_3706_), .B(_3704_), .C(raddr1_2_bF_buf7_), .Y(_3707_) );
OAI21X1 OAI21X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_1458_), .B(raddr1_0_bF_buf5_), .C(raddr1_1_bF_buf11_bF_buf2_), .Y(_3708_) );
AOI21X1 AOI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(regs_20__25_), .B(raddr1_0_bF_buf4_), .C(_3708_), .Y(_3709_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(regs_22__25_), .B(raddr1_0_bF_buf3_), .Y(_3710_) );
OAI21X1 OAI21X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_1360_), .B(raddr1_0_bF_buf2_), .C(_2415__bF_buf7), .Y(_3711_) );
OAI21X1 OAI21X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_3711_), .B(_3710_), .C(_2399__bF_buf2), .Y(_3712_) );
OAI22X1 OAI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_3703_), .B(_3707_), .C(_3712_), .D(_3709_), .Y(_3713_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(regs_29__25_), .Y(_3714_) );
NAND2X1 NAND2X1_618 ( .gnd(gnd), .vdd(vdd), .A(regs_28__25_), .B(raddr1_0_bF_buf1_), .Y(_3715_) );
OAI21X1 OAI21X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_3714_), .B(raddr1_0_bF_buf0_), .C(_3715_), .Y(_3716_) );
MUX2X1 MUX2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_3716_), .B(regs_30__25_), .S(raddr1_1_bF_buf10_bF_buf2_), .Y(_3717_) );
NAND2X1 NAND2X1_619 ( .gnd(gnd), .vdd(vdd), .A(regs_26__25_), .B(raddr1_0_bF_buf96_), .Y(_3718_) );
OAI21X1 OAI21X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_1193_), .B(raddr1_0_bF_buf95_), .C(_3718_), .Y(_3719_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(regs_25__25_), .Y(_3720_) );
NAND2X1 NAND2X1_620 ( .gnd(gnd), .vdd(vdd), .A(regs_24__25_), .B(raddr1_0_bF_buf94_), .Y(_3721_) );
OAI21X1 OAI21X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_3720_), .B(raddr1_0_bF_buf93_), .C(_3721_), .Y(_3722_) );
MUX2X1 MUX2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_3722_), .B(_3719_), .S(raddr1_1_bF_buf9_bF_buf2_), .Y(_3723_) );
MUX2X1 MUX2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_3723_), .B(_3717_), .S(raddr1_2_bF_buf6_), .Y(_3724_) );
MUX2X1 MUX2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_3724_), .B(_3713_), .S(_2398__bF_buf3), .Y(_3725_) );
MUX2X1 MUX2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_3701_), .B(_3725_), .S(raddr1_4_bF_buf4_), .Y(_5511__25_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(regs_5__26_), .Y(_3726_) );
OAI21X1 OAI21X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_3726_), .B(raddr1_0_bF_buf92_), .C(raddr1_1_bF_buf8_), .Y(_3727_) );
AOI21X1 AOI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(regs_4__26_), .B(raddr1_0_bF_buf91_), .C(_3727_), .Y(_3728_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(regs_6__26_), .B(raddr1_0_bF_buf90_), .Y(_3729_) );
OAI21X1 OAI21X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_2153_), .B(raddr1_0_bF_buf89_), .C(_2415__bF_buf6), .Y(_3730_) );
OAI21X1 OAI21X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_3730_), .B(_3729_), .C(_2399__bF_buf1), .Y(_3731_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(regs_1__26_), .Y(_3732_) );
OAI21X1 OAI21X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_3732_), .B(raddr1_0_bF_buf88_), .C(raddr1_1_bF_buf7_), .Y(_3733_) );
AOI21X1 AOI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(regs_0__26_), .B(raddr1_0_bF_buf87_), .C(_3733_), .Y(_3734_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(regs_3__26_), .Y(_3735_) );
NOR2X1 NOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf86_), .B(_3735_), .Y(_3736_) );
NAND2X1 NAND2X1_621 ( .gnd(gnd), .vdd(vdd), .A(regs_2__26_), .B(raddr1_0_bF_buf85_), .Y(_3737_) );
NAND2X1 NAND2X1_622 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf5), .B(_3737_), .Y(_3738_) );
OAI21X1 OAI21X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_3738_), .B(_3736_), .C(raddr1_2_bF_buf5_), .Y(_3739_) );
OAI22X1 OAI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(_3734_), .B(_3739_), .C(_3731_), .D(_3728_), .Y(_3740_) );
NAND2X1 NAND2X1_623 ( .gnd(gnd), .vdd(vdd), .A(regs_10__26_), .B(raddr1_0_bF_buf84_), .Y(_3741_) );
OAI21X1 OAI21X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_1954_), .B(raddr1_0_bF_buf83_), .C(_3741_), .Y(_3742_) );
NAND2X1 NAND2X1_624 ( .gnd(gnd), .vdd(vdd), .A(regs_8__26_), .B(raddr1_0_bF_buf82_), .Y(_3743_) );
OAI21X1 OAI21X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_2052_), .B(raddr1_0_bF_buf81_), .C(_3743_), .Y(_3744_) );
MUX2X1 MUX2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_3744_), .B(_3742_), .S(raddr1_1_bF_buf6_), .Y(_3745_) );
NAND2X1 NAND2X1_625 ( .gnd(gnd), .vdd(vdd), .A(regs_14__26_), .B(raddr1_0_bF_buf80_), .Y(_3746_) );
OAI21X1 OAI21X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_1757_), .B(raddr1_0_bF_buf79_), .C(_3746_), .Y(_3747_) );
NAND2X1 NAND2X1_626 ( .gnd(gnd), .vdd(vdd), .A(regs_12__26_), .B(raddr1_0_bF_buf78_), .Y(_3748_) );
OAI21X1 OAI21X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_1855_), .B(raddr1_0_bF_buf77_), .C(_3748_), .Y(_3749_) );
MUX2X1 MUX2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_3749_), .B(_3747_), .S(raddr1_1_bF_buf5_), .Y(_3750_) );
MUX2X1 MUX2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_3750_), .B(_3745_), .S(_2399__bF_buf0), .Y(_3751_) );
MUX2X1 MUX2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_3751_), .B(_3740_), .S(_2398__bF_buf2), .Y(_3752_) );
OAI21X1 OAI21X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_1657_), .B(raddr1_0_bF_buf76_), .C(raddr1_1_bF_buf4_), .Y(_3753_) );
AOI21X1 AOI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(regs_16__26_), .B(raddr1_0_bF_buf75_), .C(_3753_), .Y(_3754_) );
NOR2X1 NOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf74_), .B(_1559_), .Y(_3755_) );
NAND2X1 NAND2X1_627 ( .gnd(gnd), .vdd(vdd), .A(regs_18__26_), .B(raddr1_0_bF_buf73_), .Y(_3756_) );
NAND2X1 NAND2X1_628 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf4), .B(_3756_), .Y(_3757_) );
OAI21X1 OAI21X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_3757_), .B(_3755_), .C(raddr1_2_bF_buf4_), .Y(_3758_) );
OAI21X1 OAI21X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_1460_), .B(raddr1_0_bF_buf72_), .C(raddr1_1_bF_buf3_), .Y(_3759_) );
AOI21X1 AOI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(regs_20__26_), .B(raddr1_0_bF_buf71_), .C(_3759_), .Y(_3760_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(regs_22__26_), .B(raddr1_0_bF_buf70_), .Y(_3761_) );
OAI21X1 OAI21X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_1362_), .B(raddr1_0_bF_buf69_), .C(_2415__bF_buf3), .Y(_3762_) );
OAI21X1 OAI21X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_3762_), .B(_3761_), .C(_2399__bF_buf8), .Y(_3763_) );
OAI22X1 OAI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_3754_), .B(_3758_), .C(_3763_), .D(_3760_), .Y(_3764_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(regs_29__26_), .Y(_3765_) );
NAND2X1 NAND2X1_629 ( .gnd(gnd), .vdd(vdd), .A(regs_28__26_), .B(raddr1_0_bF_buf68_), .Y(_3766_) );
OAI21X1 OAI21X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_3765_), .B(raddr1_0_bF_buf67_), .C(_3766_), .Y(_3767_) );
MUX2X1 MUX2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_3767_), .B(regs_30__26_), .S(raddr1_1_bF_buf2_), .Y(_3768_) );
NAND2X1 NAND2X1_630 ( .gnd(gnd), .vdd(vdd), .A(regs_26__26_), .B(raddr1_0_bF_buf66_), .Y(_3769_) );
OAI21X1 OAI21X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(raddr1_0_bF_buf65_), .C(_3769_), .Y(_3770_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(regs_25__26_), .Y(_3771_) );
NAND2X1 NAND2X1_631 ( .gnd(gnd), .vdd(vdd), .A(regs_24__26_), .B(raddr1_0_bF_buf64_), .Y(_3772_) );
OAI21X1 OAI21X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_3771_), .B(raddr1_0_bF_buf63_), .C(_3772_), .Y(_3773_) );
MUX2X1 MUX2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_3773_), .B(_3770_), .S(raddr1_1_bF_buf1_), .Y(_3774_) );
MUX2X1 MUX2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_3774_), .B(_3768_), .S(raddr1_2_bF_buf3_), .Y(_3775_) );
MUX2X1 MUX2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_3775_), .B(_3764_), .S(_2398__bF_buf1), .Y(_3776_) );
MUX2X1 MUX2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_3752_), .B(_3776_), .S(raddr1_4_bF_buf3_), .Y(_5511__26_) );
NAND2X1 NAND2X1_632 ( .gnd(gnd), .vdd(vdd), .A(regs_22__27_), .B(raddr1_0_bF_buf62_), .Y(_3777_) );
OAI21X1 OAI21X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_1364_), .B(raddr1_0_bF_buf61_), .C(_3777_), .Y(_3778_) );
NAND2X1 NAND2X1_633 ( .gnd(gnd), .vdd(vdd), .A(regs_20__27_), .B(raddr1_0_bF_buf60_), .Y(_3779_) );
OAI21X1 OAI21X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_1462_), .B(raddr1_0_bF_buf59_), .C(_3779_), .Y(_3780_) );
MUX2X1 MUX2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_3780_), .B(_3778_), .S(raddr1_1_bF_buf0_), .Y(_3781_) );
NAND2X1 NAND2X1_634 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf7), .B(_3781_), .Y(_3782_) );
NAND2X1 NAND2X1_635 ( .gnd(gnd), .vdd(vdd), .A(regs_18__27_), .B(raddr1_0_bF_buf58_), .Y(_3783_) );
OAI21X1 OAI21X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .B(raddr1_0_bF_buf57_), .C(_3783_), .Y(_3784_) );
NAND2X1 NAND2X1_636 ( .gnd(gnd), .vdd(vdd), .A(regs_16__27_), .B(raddr1_0_bF_buf56_), .Y(_3785_) );
OAI21X1 OAI21X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_1659_), .B(raddr1_0_bF_buf55_), .C(_3785_), .Y(_3786_) );
MUX2X1 MUX2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_3786_), .B(_3784_), .S(raddr1_1_bF_buf14_bF_buf1_), .Y(_3787_) );
AOI21X1 AOI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(raddr1_2_bF_buf2_), .B(_3787_), .C(_2398__bF_buf0), .Y(_3788_) );
OAI21X1 OAI21X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(raddr1_0_bF_buf54_), .C(raddr1_2_bF_buf1_), .Y(_3789_) );
AOI21X1 AOI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(regs_26__27_), .B(raddr1_0_bF_buf53_), .C(_3789_), .Y(_3790_) );
OAI21X1 OAI21X1_1503 ( .gnd(gnd), .vdd(vdd), .A(regs_30__27_), .B(raddr1_2_bF_buf0_), .C(_2415__bF_buf2), .Y(_3791_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(regs_25__27_), .Y(_3792_) );
OAI21X1 OAI21X1_1504 ( .gnd(gnd), .vdd(vdd), .A(_3792_), .B(raddr1_0_bF_buf52_), .C(raddr1_2_bF_buf10_), .Y(_3793_) );
AOI21X1 AOI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(regs_24__27_), .B(raddr1_0_bF_buf51_), .C(_3793_), .Y(_3794_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(regs_29__27_), .Y(_3795_) );
NOR2X1 NOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf50_), .B(_3795_), .Y(_3796_) );
NAND2X1 NAND2X1_637 ( .gnd(gnd), .vdd(vdd), .A(regs_28__27_), .B(raddr1_0_bF_buf49_), .Y(_3797_) );
NAND2X1 NAND2X1_638 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf6), .B(_3797_), .Y(_3798_) );
OAI21X1 OAI21X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_3798_), .B(_3796_), .C(raddr1_1_bF_buf13_bF_buf1_), .Y(_3799_) );
OAI22X1 OAI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(_3790_), .B(_3791_), .C(_3799_), .D(_3794_), .Y(_3800_) );
AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_3800_), .B(_2398__bF_buf7), .C(_3782_), .D(_3788_), .Y(_3801_) );
NAND2X1 NAND2X1_639 ( .gnd(gnd), .vdd(vdd), .A(regs_6__27_), .B(raddr1_0_bF_buf48_), .Y(_3802_) );
OAI21X1 OAI21X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_2155_), .B(raddr1_0_bF_buf47_), .C(_3802_), .Y(_3803_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(regs_5__27_), .Y(_3804_) );
NAND2X1 NAND2X1_640 ( .gnd(gnd), .vdd(vdd), .A(regs_4__27_), .B(raddr1_0_bF_buf46_), .Y(_3805_) );
OAI21X1 OAI21X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_3804_), .B(raddr1_0_bF_buf45_), .C(_3805_), .Y(_3806_) );
MUX2X1 MUX2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_3806_), .B(_3803_), .S(raddr1_1_bF_buf12_bF_buf1_), .Y(_3807_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(regs_3__27_), .Y(_3808_) );
NAND2X1 NAND2X1_641 ( .gnd(gnd), .vdd(vdd), .A(regs_2__27_), .B(raddr1_0_bF_buf44_), .Y(_3809_) );
OAI21X1 OAI21X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_3808_), .B(raddr1_0_bF_buf43_), .C(_3809_), .Y(_3810_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(regs_1__27_), .Y(_3811_) );
NAND2X1 NAND2X1_642 ( .gnd(gnd), .vdd(vdd), .A(regs_0__27_), .B(raddr1_0_bF_buf42_), .Y(_3812_) );
OAI21X1 OAI21X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_3811_), .B(raddr1_0_bF_buf41_), .C(_3812_), .Y(_3813_) );
MUX2X1 MUX2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_3813_), .B(_3810_), .S(raddr1_1_bF_buf11_bF_buf1_), .Y(_3814_) );
MUX2X1 MUX2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_3814_), .B(_3807_), .S(raddr1_2_bF_buf9_), .Y(_3815_) );
NAND2X1 NAND2X1_643 ( .gnd(gnd), .vdd(vdd), .A(regs_14__27_), .B(raddr1_0_bF_buf40_), .Y(_3816_) );
OAI21X1 OAI21X1_1510 ( .gnd(gnd), .vdd(vdd), .A(_1759_), .B(raddr1_0_bF_buf39_), .C(_3816_), .Y(_3817_) );
NAND2X1 NAND2X1_644 ( .gnd(gnd), .vdd(vdd), .A(regs_12__27_), .B(raddr1_0_bF_buf38_), .Y(_3818_) );
OAI21X1 OAI21X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_1857_), .B(raddr1_0_bF_buf37_), .C(_3818_), .Y(_3819_) );
MUX2X1 MUX2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_3819_), .B(_3817_), .S(raddr1_1_bF_buf10_bF_buf1_), .Y(_3820_) );
NAND2X1 NAND2X1_645 ( .gnd(gnd), .vdd(vdd), .A(regs_10__27_), .B(raddr1_0_bF_buf36_), .Y(_3821_) );
OAI21X1 OAI21X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_1956_), .B(raddr1_0_bF_buf35_), .C(_3821_), .Y(_3822_) );
NAND2X1 NAND2X1_646 ( .gnd(gnd), .vdd(vdd), .A(regs_8__27_), .B(raddr1_0_bF_buf34_), .Y(_3823_) );
OAI21X1 OAI21X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_2054_), .B(raddr1_0_bF_buf33_), .C(_3823_), .Y(_3824_) );
MUX2X1 MUX2X1_262 ( .gnd(gnd), .vdd(vdd), .A(_3824_), .B(_3822_), .S(raddr1_1_bF_buf9_bF_buf1_), .Y(_3825_) );
MUX2X1 MUX2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_3825_), .B(_3820_), .S(raddr1_2_bF_buf8_), .Y(_3826_) );
MUX2X1 MUX2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_3826_), .B(_3815_), .S(_2398__bF_buf6), .Y(_3827_) );
MUX2X1 MUX2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_3827_), .B(_3801_), .S(raddr1_4_bF_buf2_), .Y(_5511__27_) );
NAND2X1 NAND2X1_647 ( .gnd(gnd), .vdd(vdd), .A(regs_22__28_), .B(raddr1_0_bF_buf32_), .Y(_3828_) );
OAI21X1 OAI21X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_1366_), .B(raddr1_0_bF_buf31_), .C(_3828_), .Y(_3829_) );
NAND2X1 NAND2X1_648 ( .gnd(gnd), .vdd(vdd), .A(regs_20__28_), .B(raddr1_0_bF_buf30_), .Y(_3830_) );
OAI21X1 OAI21X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(raddr1_0_bF_buf29_), .C(_3830_), .Y(_3831_) );
MUX2X1 MUX2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_3831_), .B(_3829_), .S(raddr1_1_bF_buf8_), .Y(_3832_) );
NAND2X1 NAND2X1_649 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf5), .B(_3832_), .Y(_3833_) );
NAND2X1 NAND2X1_650 ( .gnd(gnd), .vdd(vdd), .A(regs_18__28_), .B(raddr1_0_bF_buf28_), .Y(_3834_) );
OAI21X1 OAI21X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_1563_), .B(raddr1_0_bF_buf27_), .C(_3834_), .Y(_3835_) );
NAND2X1 NAND2X1_651 ( .gnd(gnd), .vdd(vdd), .A(regs_16__28_), .B(raddr1_0_bF_buf26_), .Y(_3836_) );
OAI21X1 OAI21X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_1661_), .B(raddr1_0_bF_buf25_), .C(_3836_), .Y(_3837_) );
MUX2X1 MUX2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_3837_), .B(_3835_), .S(raddr1_1_bF_buf7_), .Y(_3838_) );
AOI21X1 AOI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(raddr1_2_bF_buf7_), .B(_3838_), .C(_2398__bF_buf5), .Y(_3839_) );
OAI21X1 OAI21X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_1199_), .B(raddr1_0_bF_buf24_), .C(raddr1_2_bF_buf6_), .Y(_3840_) );
AOI21X1 AOI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(regs_26__28_), .B(raddr1_0_bF_buf23_), .C(_3840_), .Y(_3841_) );
OAI21X1 OAI21X1_1519 ( .gnd(gnd), .vdd(vdd), .A(regs_30__28_), .B(raddr1_2_bF_buf5_), .C(_2415__bF_buf1), .Y(_3842_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(regs_25__28_), .Y(_3843_) );
OAI21X1 OAI21X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_3843_), .B(raddr1_0_bF_buf22_), .C(raddr1_2_bF_buf4_), .Y(_3844_) );
AOI21X1 AOI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(regs_24__28_), .B(raddr1_0_bF_buf21_), .C(_3844_), .Y(_3845_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(regs_29__28_), .Y(_3846_) );
NOR2X1 NOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf20_), .B(_3846_), .Y(_3847_) );
NAND2X1 NAND2X1_652 ( .gnd(gnd), .vdd(vdd), .A(regs_28__28_), .B(raddr1_0_bF_buf19_), .Y(_3848_) );
NAND2X1 NAND2X1_653 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf4), .B(_3848_), .Y(_3849_) );
OAI21X1 OAI21X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_3849_), .B(_3847_), .C(raddr1_1_bF_buf6_), .Y(_3850_) );
OAI22X1 OAI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_3841_), .B(_3842_), .C(_3850_), .D(_3845_), .Y(_3851_) );
AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_3851_), .B(_2398__bF_buf4), .C(_3833_), .D(_3839_), .Y(_3852_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(regs_5__28_), .Y(_3853_) );
OAI21X1 OAI21X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_3853_), .B(raddr1_0_bF_buf18_), .C(raddr1_1_bF_buf5_), .Y(_3854_) );
AOI21X1 AOI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(regs_4__28_), .B(raddr1_0_bF_buf17_), .C(_3854_), .Y(_3855_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(regs_6__28_), .B(raddr1_0_bF_buf16_), .Y(_3856_) );
OAI21X1 OAI21X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_2157_), .B(raddr1_0_bF_buf15_), .C(_2415__bF_buf0), .Y(_3857_) );
OAI21X1 OAI21X1_1524 ( .gnd(gnd), .vdd(vdd), .A(_3857_), .B(_3856_), .C(_2399__bF_buf3), .Y(_3858_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(regs_1__28_), .Y(_3859_) );
OAI21X1 OAI21X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_3859_), .B(raddr1_0_bF_buf14_), .C(raddr1_1_bF_buf4_), .Y(_3860_) );
AOI21X1 AOI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(regs_0__28_), .B(raddr1_0_bF_buf13_), .C(_3860_), .Y(_3861_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(regs_3__28_), .Y(_3862_) );
NOR2X1 NOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf12_), .B(_3862_), .Y(_3863_) );
NAND2X1 NAND2X1_654 ( .gnd(gnd), .vdd(vdd), .A(regs_2__28_), .B(raddr1_0_bF_buf11_), .Y(_3864_) );
NAND2X1 NAND2X1_655 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf8), .B(_3864_), .Y(_3865_) );
OAI21X1 OAI21X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_3865_), .B(_3863_), .C(raddr1_2_bF_buf3_), .Y(_3866_) );
OAI22X1 OAI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(_3861_), .B(_3866_), .C(_3858_), .D(_3855_), .Y(_3867_) );
NAND2X1 NAND2X1_656 ( .gnd(gnd), .vdd(vdd), .A(regs_10__28_), .B(raddr1_0_bF_buf10_), .Y(_3868_) );
OAI21X1 OAI21X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_1958_), .B(raddr1_0_bF_buf9_), .C(_3868_), .Y(_3869_) );
NAND2X1 NAND2X1_657 ( .gnd(gnd), .vdd(vdd), .A(regs_8__28_), .B(raddr1_0_bF_buf8_), .Y(_3870_) );
OAI21X1 OAI21X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_2056_), .B(raddr1_0_bF_buf7_), .C(_3870_), .Y(_3871_) );
MUX2X1 MUX2X1_268 ( .gnd(gnd), .vdd(vdd), .A(_3871_), .B(_3869_), .S(raddr1_1_bF_buf3_), .Y(_3872_) );
NAND2X1 NAND2X1_658 ( .gnd(gnd), .vdd(vdd), .A(regs_14__28_), .B(raddr1_0_bF_buf6_), .Y(_3873_) );
OAI21X1 OAI21X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_1761_), .B(raddr1_0_bF_buf5_), .C(_3873_), .Y(_3874_) );
NAND2X1 NAND2X1_659 ( .gnd(gnd), .vdd(vdd), .A(regs_12__28_), .B(raddr1_0_bF_buf4_), .Y(_3875_) );
OAI21X1 OAI21X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_1859_), .B(raddr1_0_bF_buf3_), .C(_3875_), .Y(_3876_) );
MUX2X1 MUX2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_3876_), .B(_3874_), .S(raddr1_1_bF_buf2_), .Y(_3877_) );
MUX2X1 MUX2X1_270 ( .gnd(gnd), .vdd(vdd), .A(_3877_), .B(_3872_), .S(_2399__bF_buf2), .Y(_3878_) );
MUX2X1 MUX2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_3878_), .B(_3867_), .S(_2398__bF_buf3), .Y(_3879_) );
MUX2X1 MUX2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_3879_), .B(_3852_), .S(raddr1_4_bF_buf1_), .Y(_5511__28_) );
NAND2X1 NAND2X1_660 ( .gnd(gnd), .vdd(vdd), .A(regs_22__29_), .B(raddr1_0_bF_buf2_), .Y(_3880_) );
OAI21X1 OAI21X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_1368_), .B(raddr1_0_bF_buf1_), .C(_3880_), .Y(_3881_) );
NAND2X1 NAND2X1_661 ( .gnd(gnd), .vdd(vdd), .A(regs_20__29_), .B(raddr1_0_bF_buf0_), .Y(_3882_) );
OAI21X1 OAI21X1_1532 ( .gnd(gnd), .vdd(vdd), .A(_1466_), .B(raddr1_0_bF_buf96_), .C(_3882_), .Y(_3883_) );
MUX2X1 MUX2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_3883_), .B(_3881_), .S(raddr1_1_bF_buf1_), .Y(_3884_) );
NAND2X1 NAND2X1_662 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf1), .B(_3884_), .Y(_3885_) );
NAND2X1 NAND2X1_663 ( .gnd(gnd), .vdd(vdd), .A(regs_18__29_), .B(raddr1_0_bF_buf95_), .Y(_3886_) );
OAI21X1 OAI21X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_1565_), .B(raddr1_0_bF_buf94_), .C(_3886_), .Y(_3887_) );
NAND2X1 NAND2X1_664 ( .gnd(gnd), .vdd(vdd), .A(regs_16__29_), .B(raddr1_0_bF_buf93_), .Y(_3888_) );
OAI21X1 OAI21X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_1663_), .B(raddr1_0_bF_buf92_), .C(_3888_), .Y(_3889_) );
MUX2X1 MUX2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_3889_), .B(_3887_), .S(raddr1_1_bF_buf0_), .Y(_3890_) );
AOI21X1 AOI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(raddr1_2_bF_buf2_), .B(_3890_), .C(_2398__bF_buf2), .Y(_3891_) );
OAI21X1 OAI21X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_1201_), .B(raddr1_0_bF_buf91_), .C(raddr1_2_bF_buf1_), .Y(_3892_) );
AOI21X1 AOI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(regs_26__29_), .B(raddr1_0_bF_buf90_), .C(_3892_), .Y(_3893_) );
OAI21X1 OAI21X1_1536 ( .gnd(gnd), .vdd(vdd), .A(regs_30__29_), .B(raddr1_2_bF_buf0_), .C(_2415__bF_buf7), .Y(_3894_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(regs_25__29_), .Y(_3895_) );
OAI21X1 OAI21X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_3895_), .B(raddr1_0_bF_buf89_), .C(raddr1_2_bF_buf10_), .Y(_3896_) );
AOI21X1 AOI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(regs_24__29_), .B(raddr1_0_bF_buf88_), .C(_3896_), .Y(_3897_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(regs_29__29_), .Y(_3898_) );
NOR2X1 NOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf87_), .B(_3898_), .Y(_3899_) );
NAND2X1 NAND2X1_665 ( .gnd(gnd), .vdd(vdd), .A(regs_28__29_), .B(raddr1_0_bF_buf86_), .Y(_3900_) );
NAND2X1 NAND2X1_666 ( .gnd(gnd), .vdd(vdd), .A(_2399__bF_buf0), .B(_3900_), .Y(_3901_) );
OAI21X1 OAI21X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_3901_), .B(_3899_), .C(raddr1_1_bF_buf14_bF_buf0_), .Y(_3902_) );
OAI22X1 OAI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(_3893_), .B(_3894_), .C(_3902_), .D(_3897_), .Y(_3903_) );
AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_3903_), .B(_2398__bF_buf1), .C(_3885_), .D(_3891_), .Y(_3904_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(regs_5__29_), .Y(_3905_) );
OAI21X1 OAI21X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_3905_), .B(raddr1_0_bF_buf85_), .C(raddr1_1_bF_buf13_bF_buf0_), .Y(_3906_) );
AOI21X1 AOI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(regs_4__29_), .B(raddr1_0_bF_buf84_), .C(_3906_), .Y(_3907_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(regs_6__29_), .B(raddr1_0_bF_buf83_), .Y(_3908_) );
OAI21X1 OAI21X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_2159_), .B(raddr1_0_bF_buf82_), .C(_2415__bF_buf6), .Y(_3909_) );
OAI21X1 OAI21X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_3909_), .B(_3908_), .C(_2399__bF_buf8), .Y(_3910_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(regs_1__29_), .Y(_3911_) );
OAI21X1 OAI21X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_3911_), .B(raddr1_0_bF_buf81_), .C(raddr1_1_bF_buf12_bF_buf0_), .Y(_3912_) );
AOI21X1 AOI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(regs_0__29_), .B(raddr1_0_bF_buf80_), .C(_3912_), .Y(_3913_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(regs_3__29_), .Y(_3914_) );
NOR2X1 NOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf79_), .B(_3914_), .Y(_3915_) );
NAND2X1 NAND2X1_667 ( .gnd(gnd), .vdd(vdd), .A(regs_2__29_), .B(raddr1_0_bF_buf78_), .Y(_3916_) );
NAND2X1 NAND2X1_668 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf5), .B(_3916_), .Y(_3917_) );
OAI21X1 OAI21X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_3917_), .B(_3915_), .C(raddr1_2_bF_buf9_), .Y(_3918_) );
OAI22X1 OAI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(_3913_), .B(_3918_), .C(_3910_), .D(_3907_), .Y(_3919_) );
NAND2X1 NAND2X1_669 ( .gnd(gnd), .vdd(vdd), .A(regs_10__29_), .B(raddr1_0_bF_buf77_), .Y(_3920_) );
OAI21X1 OAI21X1_1544 ( .gnd(gnd), .vdd(vdd), .A(_1960_), .B(raddr1_0_bF_buf76_), .C(_3920_), .Y(_3921_) );
NAND2X1 NAND2X1_670 ( .gnd(gnd), .vdd(vdd), .A(regs_8__29_), .B(raddr1_0_bF_buf75_), .Y(_3922_) );
OAI21X1 OAI21X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_2058_), .B(raddr1_0_bF_buf74_), .C(_3922_), .Y(_3923_) );
MUX2X1 MUX2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_3923_), .B(_3921_), .S(raddr1_1_bF_buf11_bF_buf0_), .Y(_3924_) );
NAND2X1 NAND2X1_671 ( .gnd(gnd), .vdd(vdd), .A(regs_14__29_), .B(raddr1_0_bF_buf73_), .Y(_3925_) );
OAI21X1 OAI21X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_1763_), .B(raddr1_0_bF_buf72_), .C(_3925_), .Y(_3926_) );
NAND2X1 NAND2X1_672 ( .gnd(gnd), .vdd(vdd), .A(regs_12__29_), .B(raddr1_0_bF_buf71_), .Y(_3927_) );
OAI21X1 OAI21X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_1861_), .B(raddr1_0_bF_buf70_), .C(_3927_), .Y(_3928_) );
MUX2X1 MUX2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_3928_), .B(_3926_), .S(raddr1_1_bF_buf10_bF_buf0_), .Y(_3929_) );
MUX2X1 MUX2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_3929_), .B(_3924_), .S(_2399__bF_buf7), .Y(_3930_) );
MUX2X1 MUX2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_3930_), .B(_3919_), .S(_2398__bF_buf0), .Y(_3931_) );
MUX2X1 MUX2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_3931_), .B(_3904_), .S(raddr1_4_bF_buf0_), .Y(_5511__29_) );
OAI21X1 OAI21X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_1468_), .B(raddr1_0_bF_buf69_), .C(raddr1_1_bF_buf9_bF_buf0_), .Y(_3932_) );
AOI21X1 AOI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(regs_20__30_), .B(raddr1_0_bF_buf68_), .C(_3932_), .Y(_3933_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(regs_22__30_), .B(raddr1_0_bF_buf67_), .Y(_3934_) );
OAI21X1 OAI21X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_1370_), .B(raddr1_0_bF_buf66_), .C(_2415__bF_buf4), .Y(_3935_) );
OAI21X1 OAI21X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_3935_), .B(_3934_), .C(_2399__bF_buf6), .Y(_3936_) );
OAI21X1 OAI21X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_1665_), .B(raddr1_0_bF_buf65_), .C(raddr1_1_bF_buf8_), .Y(_3937_) );
AOI21X1 AOI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(regs_16__30_), .B(raddr1_0_bF_buf64_), .C(_3937_), .Y(_3938_) );
NOR2X1 NOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf63_), .B(_1567_), .Y(_3939_) );
NAND2X1 NAND2X1_673 ( .gnd(gnd), .vdd(vdd), .A(regs_18__30_), .B(raddr1_0_bF_buf62_), .Y(_3940_) );
NAND2X1 NAND2X1_674 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf3), .B(_3940_), .Y(_3941_) );
OAI21X1 OAI21X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_3941_), .B(_3939_), .C(raddr1_2_bF_buf8_), .Y(_3942_) );
OAI22X1 OAI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(_3938_), .B(_3942_), .C(_3936_), .D(_3933_), .Y(_3943_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(regs_29__30_), .Y(_3944_) );
NAND2X1 NAND2X1_675 ( .gnd(gnd), .vdd(vdd), .A(regs_28__30_), .B(raddr1_0_bF_buf61_), .Y(_3945_) );
OAI21X1 OAI21X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_3944_), .B(raddr1_0_bF_buf60_), .C(_3945_), .Y(_3946_) );
MUX2X1 MUX2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_3946_), .B(regs_30__30_), .S(raddr1_1_bF_buf7_), .Y(_3947_) );
NAND2X1 NAND2X1_676 ( .gnd(gnd), .vdd(vdd), .A(regs_26__30_), .B(raddr1_0_bF_buf59_), .Y(_3948_) );
OAI21X1 OAI21X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_1203_), .B(raddr1_0_bF_buf58_), .C(_3948_), .Y(_3949_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(regs_25__30_), .Y(_3950_) );
NAND2X1 NAND2X1_677 ( .gnd(gnd), .vdd(vdd), .A(regs_24__30_), .B(raddr1_0_bF_buf57_), .Y(_3951_) );
OAI21X1 OAI21X1_1555 ( .gnd(gnd), .vdd(vdd), .A(_3950_), .B(raddr1_0_bF_buf56_), .C(_3951_), .Y(_3952_) );
MUX2X1 MUX2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_3952_), .B(_3949_), .S(raddr1_1_bF_buf6_), .Y(_3953_) );
MUX2X1 MUX2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_3953_), .B(_3947_), .S(raddr1_2_bF_buf7_), .Y(_3954_) );
MUX2X1 MUX2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_3954_), .B(_3943_), .S(_2398__bF_buf7), .Y(_3955_) );
NAND2X1 NAND2X1_678 ( .gnd(gnd), .vdd(vdd), .A(regs_6__30_), .B(raddr1_0_bF_buf55_), .Y(_3956_) );
OAI21X1 OAI21X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_2161_), .B(raddr1_0_bF_buf54_), .C(_3956_), .Y(_3957_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(regs_5__30_), .Y(_3958_) );
NAND2X1 NAND2X1_679 ( .gnd(gnd), .vdd(vdd), .A(regs_4__30_), .B(raddr1_0_bF_buf53_), .Y(_3959_) );
OAI21X1 OAI21X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_3958_), .B(raddr1_0_bF_buf52_), .C(_3959_), .Y(_3960_) );
MUX2X1 MUX2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_3960_), .B(_3957_), .S(raddr1_1_bF_buf5_), .Y(_3961_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(regs_3__30_), .Y(_3962_) );
NAND2X1 NAND2X1_680 ( .gnd(gnd), .vdd(vdd), .A(regs_2__30_), .B(raddr1_0_bF_buf51_), .Y(_3963_) );
OAI21X1 OAI21X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_3962_), .B(raddr1_0_bF_buf50_), .C(_3963_), .Y(_3964_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(regs_1__30_), .Y(_3965_) );
NAND2X1 NAND2X1_681 ( .gnd(gnd), .vdd(vdd), .A(regs_0__30_), .B(raddr1_0_bF_buf49_), .Y(_3966_) );
OAI21X1 OAI21X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_3965_), .B(raddr1_0_bF_buf48_), .C(_3966_), .Y(_3967_) );
MUX2X1 MUX2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_3967_), .B(_3964_), .S(raddr1_1_bF_buf4_), .Y(_3968_) );
MUX2X1 MUX2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_3968_), .B(_3961_), .S(raddr1_2_bF_buf6_), .Y(_3969_) );
NAND2X1 NAND2X1_682 ( .gnd(gnd), .vdd(vdd), .A(regs_10__30_), .B(raddr1_0_bF_buf47_), .Y(_3970_) );
OAI21X1 OAI21X1_1560 ( .gnd(gnd), .vdd(vdd), .A(_1962_), .B(raddr1_0_bF_buf46_), .C(_3970_), .Y(_3971_) );
NAND2X1 NAND2X1_683 ( .gnd(gnd), .vdd(vdd), .A(regs_8__30_), .B(raddr1_0_bF_buf45_), .Y(_3972_) );
OAI21X1 OAI21X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_2060_), .B(raddr1_0_bF_buf44_), .C(_3972_), .Y(_3973_) );
MUX2X1 MUX2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_3973_), .B(_3971_), .S(raddr1_1_bF_buf3_), .Y(_3974_) );
NAND2X1 NAND2X1_684 ( .gnd(gnd), .vdd(vdd), .A(regs_14__30_), .B(raddr1_0_bF_buf43_), .Y(_3975_) );
OAI21X1 OAI21X1_1562 ( .gnd(gnd), .vdd(vdd), .A(_1765_), .B(raddr1_0_bF_buf42_), .C(_3975_), .Y(_3976_) );
NAND2X1 NAND2X1_685 ( .gnd(gnd), .vdd(vdd), .A(regs_12__30_), .B(raddr1_0_bF_buf41_), .Y(_3977_) );
OAI21X1 OAI21X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_1863_), .B(raddr1_0_bF_buf40_), .C(_3977_), .Y(_3978_) );
MUX2X1 MUX2X1_288 ( .gnd(gnd), .vdd(vdd), .A(_3978_), .B(_3976_), .S(raddr1_1_bF_buf2_), .Y(_3979_) );
MUX2X1 MUX2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_3979_), .B(_3974_), .S(_2399__bF_buf5), .Y(_3980_) );
MUX2X1 MUX2X1_290 ( .gnd(gnd), .vdd(vdd), .A(_3980_), .B(_3969_), .S(_2398__bF_buf6), .Y(_3981_) );
MUX2X1 MUX2X1_291 ( .gnd(gnd), .vdd(vdd), .A(_3981_), .B(_3955_), .S(raddr1_4_bF_buf4_), .Y(_5511__30_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(regs_5__31_), .Y(_3982_) );
OAI21X1 OAI21X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_3982_), .B(raddr1_0_bF_buf39_), .C(raddr1_1_bF_buf1_), .Y(_3983_) );
AOI21X1 AOI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(regs_4__31_), .B(raddr1_0_bF_buf38_), .C(_3983_), .Y(_3984_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(regs_6__31_), .B(raddr1_0_bF_buf37_), .Y(_3985_) );
OAI21X1 OAI21X1_1565 ( .gnd(gnd), .vdd(vdd), .A(_2163_), .B(raddr1_0_bF_buf36_), .C(_2415__bF_buf2), .Y(_3986_) );
OAI21X1 OAI21X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_3986_), .B(_3985_), .C(_2399__bF_buf4), .Y(_3987_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(regs_1__31_), .Y(_3988_) );
OAI21X1 OAI21X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_3988_), .B(raddr1_0_bF_buf35_), .C(raddr1_1_bF_buf0_), .Y(_3989_) );
AOI21X1 AOI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(regs_0__31_), .B(raddr1_0_bF_buf34_), .C(_3989_), .Y(_3990_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(regs_3__31_), .Y(_3991_) );
NOR2X1 NOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf33_), .B(_3991_), .Y(_3992_) );
NAND2X1 NAND2X1_686 ( .gnd(gnd), .vdd(vdd), .A(regs_2__31_), .B(raddr1_0_bF_buf32_), .Y(_3993_) );
NAND2X1 NAND2X1_687 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf1), .B(_3993_), .Y(_3994_) );
OAI21X1 OAI21X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_3994_), .B(_3992_), .C(raddr1_2_bF_buf5_), .Y(_3995_) );
OAI22X1 OAI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(_3990_), .B(_3995_), .C(_3987_), .D(_3984_), .Y(_3996_) );
NAND2X1 NAND2X1_688 ( .gnd(gnd), .vdd(vdd), .A(regs_10__31_), .B(raddr1_0_bF_buf31_), .Y(_3997_) );
OAI21X1 OAI21X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_1964_), .B(raddr1_0_bF_buf30_), .C(_3997_), .Y(_3998_) );
NAND2X1 NAND2X1_689 ( .gnd(gnd), .vdd(vdd), .A(regs_8__31_), .B(raddr1_0_bF_buf29_), .Y(_3999_) );
OAI21X1 OAI21X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_2062_), .B(raddr1_0_bF_buf28_), .C(_3999_), .Y(_4000_) );
MUX2X1 MUX2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_4000_), .B(_3998_), .S(raddr1_1_bF_buf14_bF_buf3_), .Y(_4001_) );
NAND2X1 NAND2X1_690 ( .gnd(gnd), .vdd(vdd), .A(regs_14__31_), .B(raddr1_0_bF_buf27_), .Y(_4002_) );
OAI21X1 OAI21X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_1767_), .B(raddr1_0_bF_buf26_), .C(_4002_), .Y(_4003_) );
NAND2X1 NAND2X1_691 ( .gnd(gnd), .vdd(vdd), .A(regs_12__31_), .B(raddr1_0_bF_buf25_), .Y(_4004_) );
OAI21X1 OAI21X1_1572 ( .gnd(gnd), .vdd(vdd), .A(_1865_), .B(raddr1_0_bF_buf24_), .C(_4004_), .Y(_4005_) );
MUX2X1 MUX2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_4005_), .B(_4003_), .S(raddr1_1_bF_buf13_bF_buf3_), .Y(_4006_) );
MUX2X1 MUX2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_4006_), .B(_4001_), .S(_2399__bF_buf3), .Y(_4007_) );
MUX2X1 MUX2X1_295 ( .gnd(gnd), .vdd(vdd), .A(_4007_), .B(_3996_), .S(_2398__bF_buf5), .Y(_4008_) );
OAI21X1 OAI21X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_1667_), .B(raddr1_0_bF_buf23_), .C(raddr1_1_bF_buf12_bF_buf3_), .Y(_4009_) );
AOI21X1 AOI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(regs_16__31_), .B(raddr1_0_bF_buf22_), .C(_4009_), .Y(_4010_) );
NOR2X1 NOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(raddr1_0_bF_buf21_), .B(_1569_), .Y(_4011_) );
NAND2X1 NAND2X1_692 ( .gnd(gnd), .vdd(vdd), .A(regs_18__31_), .B(raddr1_0_bF_buf20_), .Y(_4012_) );
NAND2X1 NAND2X1_693 ( .gnd(gnd), .vdd(vdd), .A(_2415__bF_buf0), .B(_4012_), .Y(_4013_) );
OAI21X1 OAI21X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_4013_), .B(_4011_), .C(raddr1_2_bF_buf4_), .Y(_4014_) );
OAI21X1 OAI21X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_1470_), .B(raddr1_0_bF_buf19_), .C(raddr1_1_bF_buf11_bF_buf3_), .Y(_4015_) );
AOI21X1 AOI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(regs_20__31_), .B(raddr1_0_bF_buf18_), .C(_4015_), .Y(_4016_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(regs_22__31_), .B(raddr1_0_bF_buf17_), .Y(_4017_) );
OAI21X1 OAI21X1_1576 ( .gnd(gnd), .vdd(vdd), .A(_1372_), .B(raddr1_0_bF_buf16_), .C(_2415__bF_buf8), .Y(_4018_) );
OAI21X1 OAI21X1_1577 ( .gnd(gnd), .vdd(vdd), .A(_4018_), .B(_4017_), .C(_2399__bF_buf2), .Y(_4019_) );
OAI22X1 OAI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(_4010_), .B(_4014_), .C(_4019_), .D(_4016_), .Y(_4020_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(regs_29__31_), .Y(_4021_) );
NAND2X1 NAND2X1_694 ( .gnd(gnd), .vdd(vdd), .A(regs_28__31_), .B(raddr1_0_bF_buf15_), .Y(_4022_) );
OAI21X1 OAI21X1_1578 ( .gnd(gnd), .vdd(vdd), .A(_4021_), .B(raddr1_0_bF_buf14_), .C(_4022_), .Y(_4023_) );
MUX2X1 MUX2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_4023_), .B(regs_30__31_), .S(raddr1_1_bF_buf10_bF_buf3_), .Y(_4024_) );
NAND2X1 NAND2X1_695 ( .gnd(gnd), .vdd(vdd), .A(regs_26__31_), .B(raddr1_0_bF_buf13_), .Y(_4025_) );
OAI21X1 OAI21X1_1579 ( .gnd(gnd), .vdd(vdd), .A(_1205_), .B(raddr1_0_bF_buf12_), .C(_4025_), .Y(_4026_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(regs_25__31_), .Y(_4027_) );
NAND2X1 NAND2X1_696 ( .gnd(gnd), .vdd(vdd), .A(regs_24__31_), .B(raddr1_0_bF_buf11_), .Y(_4028_) );
OAI21X1 OAI21X1_1580 ( .gnd(gnd), .vdd(vdd), .A(_4027_), .B(raddr1_0_bF_buf10_), .C(_4028_), .Y(_4029_) );
MUX2X1 MUX2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_4029_), .B(_4026_), .S(raddr1_1_bF_buf9_bF_buf3_), .Y(_4030_) );
MUX2X1 MUX2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_4030_), .B(_4024_), .S(raddr1_2_bF_buf3_), .Y(_4031_) );
MUX2X1 MUX2X1_299 ( .gnd(gnd), .vdd(vdd), .A(_4031_), .B(_4020_), .S(_2398__bF_buf4), .Y(_4032_) );
MUX2X1 MUX2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_4008_), .B(_4032_), .S(raddr1_4_bF_buf3_), .Y(_5511__31_) );
INVX8 INVX8_5 ( .gnd(gnd), .vdd(vdd), .A(raddr2[3]), .Y(_4033_) );
OAI21X1 OAI21X1_1581 ( .gnd(gnd), .vdd(vdd), .A(_2427_), .B(raddr2_0_bF_buf96_), .C(raddr2_1_bF_buf14_bF_buf3_), .Y(_4034_) );
AOI21X1 AOI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(regs_4__0_), .B(raddr2_0_bF_buf95_), .C(_4034_), .Y(_4035_) );
INVX8 INVX8_6 ( .gnd(gnd), .vdd(vdd), .A(raddr2_2_bF_buf10_), .Y(_4036_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(regs_6__0_), .B(raddr2_0_bF_buf94_), .Y(_4037_) );
INVX8 INVX8_7 ( .gnd(gnd), .vdd(vdd), .A(raddr2_1_bF_buf13_bF_buf3_), .Y(_4038_) );
OAI21X1 OAI21X1_1582 ( .gnd(gnd), .vdd(vdd), .A(_2097_), .B(raddr2_0_bF_buf93_), .C(_4038__bF_buf8), .Y(_4039_) );
OAI21X1 OAI21X1_1583 ( .gnd(gnd), .vdd(vdd), .A(_4039_), .B(_4037_), .C(_4036__bF_buf8), .Y(_4040_) );
OAI21X1 OAI21X1_1584 ( .gnd(gnd), .vdd(vdd), .A(_2433_), .B(raddr2_0_bF_buf92_), .C(raddr2_1_bF_buf12_bF_buf3_), .Y(_4041_) );
AOI21X1 AOI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(regs_0__0_), .B(raddr2_0_bF_buf91_), .C(_4041_), .Y(_4042_) );
AOI21X1 AOI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(regs_2__0_), .B(raddr2_0_bF_buf90_), .C(raddr2_1_bF_buf11_), .Y(_4043_) );
OAI21X1 OAI21X1_1585 ( .gnd(gnd), .vdd(vdd), .A(_2436_), .B(raddr2_0_bF_buf89_), .C(_4043_), .Y(_4044_) );
NAND2X1 NAND2X1_697 ( .gnd(gnd), .vdd(vdd), .A(raddr2_2_bF_buf9_), .B(_4044_), .Y(_4045_) );
OAI22X1 OAI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(_4045_), .B(_4042_), .C(_4040_), .D(_4035_), .Y(_4046_) );
NAND2X1 NAND2X1_698 ( .gnd(gnd), .vdd(vdd), .A(regs_10__0_), .B(raddr2_0_bF_buf88_), .Y(_4047_) );
OAI21X1 OAI21X1_1586 ( .gnd(gnd), .vdd(vdd), .A(_1900_), .B(raddr2_0_bF_buf87_), .C(_4047_), .Y(_4048_) );
NAND2X1 NAND2X1_699 ( .gnd(gnd), .vdd(vdd), .A(regs_8__0_), .B(raddr2_0_bF_buf86_), .Y(_4049_) );
OAI21X1 OAI21X1_1587 ( .gnd(gnd), .vdd(vdd), .A(_1999_), .B(raddr2_0_bF_buf85_), .C(_4049_), .Y(_4050_) );
MUX2X1 MUX2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_4050_), .B(_4048_), .S(raddr2_1_bF_buf10_), .Y(_4051_) );
NAND2X1 NAND2X1_700 ( .gnd(gnd), .vdd(vdd), .A(regs_14__0_), .B(raddr2_0_bF_buf84_), .Y(_4052_) );
OAI21X1 OAI21X1_1588 ( .gnd(gnd), .vdd(vdd), .A(_1702_), .B(raddr2_0_bF_buf83_), .C(_4052_), .Y(_4053_) );
NAND2X1 NAND2X1_701 ( .gnd(gnd), .vdd(vdd), .A(regs_12__0_), .B(raddr2_0_bF_buf82_), .Y(_4054_) );
OAI21X1 OAI21X1_1589 ( .gnd(gnd), .vdd(vdd), .A(_1802_), .B(raddr2_0_bF_buf81_), .C(_4054_), .Y(_4055_) );
MUX2X1 MUX2X1_302 ( .gnd(gnd), .vdd(vdd), .A(_4055_), .B(_4053_), .S(raddr2_1_bF_buf9_), .Y(_4056_) );
MUX2X1 MUX2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_4056_), .B(_4051_), .S(_4036__bF_buf7), .Y(_4057_) );
MUX2X1 MUX2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_4057_), .B(_4046_), .S(_4033__bF_buf7), .Y(_4058_) );
OAI21X1 OAI21X1_1590 ( .gnd(gnd), .vdd(vdd), .A(_1604_), .B(raddr2_0_bF_buf80_), .C(raddr2_1_bF_buf8_), .Y(_4059_) );
AOI21X1 AOI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(regs_16__0_), .B(raddr2_0_bF_buf79_), .C(_4059_), .Y(_4060_) );
NOR2X1 NOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf78_), .B(_1505_), .Y(_4061_) );
NAND2X1 NAND2X1_702 ( .gnd(gnd), .vdd(vdd), .A(regs_18__0_), .B(raddr2_0_bF_buf77_), .Y(_4062_) );
NAND2X1 NAND2X1_703 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf7), .B(_4062_), .Y(_4063_) );
OAI21X1 OAI21X1_1591 ( .gnd(gnd), .vdd(vdd), .A(_4063_), .B(_4061_), .C(raddr2_2_bF_buf8_), .Y(_4064_) );
OAI21X1 OAI21X1_1592 ( .gnd(gnd), .vdd(vdd), .A(_1407_), .B(raddr2_0_bF_buf76_), .C(raddr2_1_bF_buf7_), .Y(_4065_) );
AOI21X1 AOI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(regs_20__0_), .B(raddr2_0_bF_buf75_), .C(_4065_), .Y(_4066_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(regs_22__0_), .B(raddr2_0_bF_buf74_), .Y(_4067_) );
OAI21X1 OAI21X1_1593 ( .gnd(gnd), .vdd(vdd), .A(_1307_), .B(raddr2_0_bF_buf73_), .C(_4038__bF_buf6), .Y(_4068_) );
OAI21X1 OAI21X1_1594 ( .gnd(gnd), .vdd(vdd), .A(_4068_), .B(_4067_), .C(_4036__bF_buf6), .Y(_4069_) );
OAI22X1 OAI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(_4060_), .B(_4064_), .C(_4069_), .D(_4066_), .Y(_4070_) );
NAND2X1 NAND2X1_704 ( .gnd(gnd), .vdd(vdd), .A(regs_28__0_), .B(raddr2_0_bF_buf72_), .Y(_4071_) );
OAI21X1 OAI21X1_1595 ( .gnd(gnd), .vdd(vdd), .A(_2420_), .B(raddr2_0_bF_buf71_), .C(_4071_), .Y(_4072_) );
MUX2X1 MUX2X1_305 ( .gnd(gnd), .vdd(vdd), .A(_4072_), .B(regs_30__0_), .S(raddr2_1_bF_buf6_), .Y(_4073_) );
NAND2X1 NAND2X1_705 ( .gnd(gnd), .vdd(vdd), .A(regs_26__0_), .B(raddr2_0_bF_buf70_), .Y(_4074_) );
OAI21X1 OAI21X1_1596 ( .gnd(gnd), .vdd(vdd), .A(_1138_), .B(raddr2_0_bF_buf69_), .C(_4074_), .Y(_4075_) );
NAND2X1 NAND2X1_706 ( .gnd(gnd), .vdd(vdd), .A(regs_24__0_), .B(raddr2_0_bF_buf68_), .Y(_4076_) );
OAI21X1 OAI21X1_1597 ( .gnd(gnd), .vdd(vdd), .A(_2417_), .B(raddr2_0_bF_buf67_), .C(_4076_), .Y(_4077_) );
MUX2X1 MUX2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_4077_), .B(_4075_), .S(raddr2_1_bF_buf5_), .Y(_4078_) );
MUX2X1 MUX2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_4078_), .B(_4073_), .S(raddr2_2_bF_buf7_), .Y(_4079_) );
MUX2X1 MUX2X1_308 ( .gnd(gnd), .vdd(vdd), .A(_4079_), .B(_4070_), .S(_4033__bF_buf6), .Y(_4080_) );
MUX2X1 MUX2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_4058_), .B(_4080_), .S(raddr2_4_bF_buf4_), .Y(_5512__0_) );
OAI21X1 OAI21X1_1598 ( .gnd(gnd), .vdd(vdd), .A(_2479_), .B(raddr2_0_bF_buf66_), .C(raddr2_1_bF_buf4_), .Y(_4081_) );
AOI21X1 AOI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(regs_4__1_), .B(raddr2_0_bF_buf65_), .C(_4081_), .Y(_4082_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(regs_6__1_), .B(raddr2_0_bF_buf64_), .Y(_4083_) );
OAI21X1 OAI21X1_1599 ( .gnd(gnd), .vdd(vdd), .A(_2103_), .B(raddr2_0_bF_buf63_), .C(_4038__bF_buf5), .Y(_4084_) );
OAI21X1 OAI21X1_1600 ( .gnd(gnd), .vdd(vdd), .A(_4084_), .B(_4083_), .C(_4036__bF_buf5), .Y(_4085_) );
OAI21X1 OAI21X1_1601 ( .gnd(gnd), .vdd(vdd), .A(_2486_), .B(raddr2_0_bF_buf62_), .C(raddr2_1_bF_buf3_), .Y(_4086_) );
AOI21X1 AOI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(regs_0__1_), .B(raddr2_0_bF_buf61_), .C(_4086_), .Y(_4087_) );
NOR2X1 NOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf60_), .B(_2483_), .Y(_4088_) );
NAND2X1 NAND2X1_707 ( .gnd(gnd), .vdd(vdd), .A(regs_2__1_), .B(raddr2_0_bF_buf59_), .Y(_4089_) );
NAND2X1 NAND2X1_708 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf4), .B(_4089_), .Y(_4090_) );
OAI21X1 OAI21X1_1602 ( .gnd(gnd), .vdd(vdd), .A(_4090_), .B(_4088_), .C(raddr2_2_bF_buf6_), .Y(_4091_) );
OAI22X1 OAI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(_4087_), .B(_4091_), .C(_4085_), .D(_4082_), .Y(_4092_) );
NAND2X1 NAND2X1_709 ( .gnd(gnd), .vdd(vdd), .A(regs_10__1_), .B(raddr2_0_bF_buf58_), .Y(_4093_) );
OAI21X1 OAI21X1_1603 ( .gnd(gnd), .vdd(vdd), .A(_1904_), .B(raddr2_0_bF_buf57_), .C(_4093_), .Y(_4094_) );
NAND2X1 NAND2X1_710 ( .gnd(gnd), .vdd(vdd), .A(regs_8__1_), .B(raddr2_0_bF_buf56_), .Y(_4095_) );
OAI21X1 OAI21X1_1604 ( .gnd(gnd), .vdd(vdd), .A(_2002_), .B(raddr2_0_bF_buf55_), .C(_4095_), .Y(_4096_) );
MUX2X1 MUX2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_4096_), .B(_4094_), .S(raddr2_1_bF_buf2_), .Y(_4097_) );
NAND2X1 NAND2X1_711 ( .gnd(gnd), .vdd(vdd), .A(regs_14__1_), .B(raddr2_0_bF_buf54_), .Y(_4098_) );
OAI21X1 OAI21X1_1605 ( .gnd(gnd), .vdd(vdd), .A(_1707_), .B(raddr2_0_bF_buf53_), .C(_4098_), .Y(_4099_) );
NAND2X1 NAND2X1_712 ( .gnd(gnd), .vdd(vdd), .A(regs_12__1_), .B(raddr2_0_bF_buf52_), .Y(_4100_) );
OAI21X1 OAI21X1_1606 ( .gnd(gnd), .vdd(vdd), .A(_1805_), .B(raddr2_0_bF_buf51_), .C(_4100_), .Y(_4101_) );
MUX2X1 MUX2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_4101_), .B(_4099_), .S(raddr2_1_bF_buf1_), .Y(_4102_) );
MUX2X1 MUX2X1_312 ( .gnd(gnd), .vdd(vdd), .A(_4102_), .B(_4097_), .S(_4036__bF_buf4), .Y(_4103_) );
MUX2X1 MUX2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_4103_), .B(_4092_), .S(_4033__bF_buf5), .Y(_4104_) );
OAI21X1 OAI21X1_1607 ( .gnd(gnd), .vdd(vdd), .A(_1607_), .B(raddr2_0_bF_buf50_), .C(raddr2_1_bF_buf0_), .Y(_4105_) );
AOI21X1 AOI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(regs_16__1_), .B(raddr2_0_bF_buf49_), .C(_4105_), .Y(_4106_) );
NOR2X1 NOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf48_), .B(_1509_), .Y(_4107_) );
NAND2X1 NAND2X1_713 ( .gnd(gnd), .vdd(vdd), .A(regs_18__1_), .B(raddr2_0_bF_buf47_), .Y(_4108_) );
NAND2X1 NAND2X1_714 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf3), .B(_4108_), .Y(_4109_) );
OAI21X1 OAI21X1_1608 ( .gnd(gnd), .vdd(vdd), .A(_4109_), .B(_4107_), .C(raddr2_2_bF_buf5_), .Y(_4110_) );
OAI21X1 OAI21X1_1609 ( .gnd(gnd), .vdd(vdd), .A(_1410_), .B(raddr2_0_bF_buf46_), .C(raddr2_1_bF_buf14_bF_buf2_), .Y(_4111_) );
AOI21X1 AOI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(regs_20__1_), .B(raddr2_0_bF_buf45_), .C(_4111_), .Y(_4112_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(regs_22__1_), .B(raddr2_0_bF_buf44_), .Y(_4113_) );
OAI21X1 OAI21X1_1610 ( .gnd(gnd), .vdd(vdd), .A(_1312_), .B(raddr2_0_bF_buf43_), .C(_4038__bF_buf2), .Y(_4114_) );
OAI21X1 OAI21X1_1611 ( .gnd(gnd), .vdd(vdd), .A(_4114_), .B(_4113_), .C(_4036__bF_buf3), .Y(_4115_) );
OAI22X1 OAI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(_4106_), .B(_4110_), .C(_4115_), .D(_4112_), .Y(_4116_) );
NAND2X1 NAND2X1_715 ( .gnd(gnd), .vdd(vdd), .A(regs_28__1_), .B(raddr2_0_bF_buf42_), .Y(_4117_) );
OAI21X1 OAI21X1_1612 ( .gnd(gnd), .vdd(vdd), .A(_2465_), .B(raddr2_0_bF_buf41_), .C(_4117_), .Y(_4118_) );
MUX2X1 MUX2X1_314 ( .gnd(gnd), .vdd(vdd), .A(_4118_), .B(regs_30__1_), .S(raddr2_1_bF_buf13_bF_buf2_), .Y(_4119_) );
NAND2X1 NAND2X1_716 ( .gnd(gnd), .vdd(vdd), .A(regs_26__1_), .B(raddr2_0_bF_buf40_), .Y(_4120_) );
OAI21X1 OAI21X1_1613 ( .gnd(gnd), .vdd(vdd), .A(_1145_), .B(raddr2_0_bF_buf39_), .C(_4120_), .Y(_4121_) );
NAND2X1 NAND2X1_717 ( .gnd(gnd), .vdd(vdd), .A(regs_24__1_), .B(raddr2_0_bF_buf38_), .Y(_4122_) );
OAI21X1 OAI21X1_1614 ( .gnd(gnd), .vdd(vdd), .A(_2471_), .B(raddr2_0_bF_buf37_), .C(_4122_), .Y(_4123_) );
MUX2X1 MUX2X1_315 ( .gnd(gnd), .vdd(vdd), .A(_4123_), .B(_4121_), .S(raddr2_1_bF_buf12_bF_buf2_), .Y(_4124_) );
MUX2X1 MUX2X1_316 ( .gnd(gnd), .vdd(vdd), .A(_4124_), .B(_4119_), .S(raddr2_2_bF_buf4_), .Y(_4125_) );
MUX2X1 MUX2X1_317 ( .gnd(gnd), .vdd(vdd), .A(_4125_), .B(_4116_), .S(_4033__bF_buf4), .Y(_4126_) );
MUX2X1 MUX2X1_318 ( .gnd(gnd), .vdd(vdd), .A(_4104_), .B(_4126_), .S(raddr2_4_bF_buf3_), .Y(_5512__1_) );
NAND2X1 NAND2X1_718 ( .gnd(gnd), .vdd(vdd), .A(regs_22__2_), .B(raddr2_0_bF_buf36_), .Y(_4127_) );
OAI21X1 OAI21X1_1615 ( .gnd(gnd), .vdd(vdd), .A(_1314_), .B(raddr2_0_bF_buf35_), .C(_4127_), .Y(_4128_) );
NAND2X1 NAND2X1_719 ( .gnd(gnd), .vdd(vdd), .A(regs_20__2_), .B(raddr2_0_bF_buf34_), .Y(_4129_) );
OAI21X1 OAI21X1_1616 ( .gnd(gnd), .vdd(vdd), .A(_1412_), .B(raddr2_0_bF_buf33_), .C(_4129_), .Y(_4130_) );
MUX2X1 MUX2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_4130_), .B(_4128_), .S(raddr2_1_bF_buf11_), .Y(_4131_) );
NAND2X1 NAND2X1_720 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf2), .B(_4131_), .Y(_4132_) );
NAND2X1 NAND2X1_721 ( .gnd(gnd), .vdd(vdd), .A(regs_18__2_), .B(raddr2_0_bF_buf32_), .Y(_4133_) );
OAI21X1 OAI21X1_1617 ( .gnd(gnd), .vdd(vdd), .A(_1511_), .B(raddr2_0_bF_buf31_), .C(_4133_), .Y(_4134_) );
NAND2X1 NAND2X1_722 ( .gnd(gnd), .vdd(vdd), .A(regs_16__2_), .B(raddr2_0_bF_buf30_), .Y(_4135_) );
OAI21X1 OAI21X1_1618 ( .gnd(gnd), .vdd(vdd), .A(_1609_), .B(raddr2_0_bF_buf29_), .C(_4135_), .Y(_4136_) );
MUX2X1 MUX2X1_320 ( .gnd(gnd), .vdd(vdd), .A(_4136_), .B(_4134_), .S(raddr2_1_bF_buf10_), .Y(_4137_) );
AOI21X1 AOI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(raddr2_2_bF_buf3_), .B(_4137_), .C(_4033__bF_buf3), .Y(_4138_) );
OAI21X1 OAI21X1_1619 ( .gnd(gnd), .vdd(vdd), .A(_1147_), .B(raddr2_0_bF_buf28_), .C(raddr2_2_bF_buf2_), .Y(_4139_) );
AOI21X1 AOI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(regs_26__2_), .B(raddr2_0_bF_buf27_), .C(_4139_), .Y(_4140_) );
OAI21X1 OAI21X1_1620 ( .gnd(gnd), .vdd(vdd), .A(regs_30__2_), .B(raddr2_2_bF_buf1_), .C(_4038__bF_buf1), .Y(_4141_) );
OAI21X1 OAI21X1_1621 ( .gnd(gnd), .vdd(vdd), .A(_2518_), .B(raddr2_0_bF_buf26_), .C(raddr2_2_bF_buf0_), .Y(_4142_) );
AOI21X1 AOI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(regs_24__2_), .B(raddr2_0_bF_buf25_), .C(_4142_), .Y(_4143_) );
NOR2X1 NOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf24_), .B(_2521_), .Y(_4144_) );
NAND2X1 NAND2X1_723 ( .gnd(gnd), .vdd(vdd), .A(regs_28__2_), .B(raddr2_0_bF_buf23_), .Y(_4145_) );
NAND2X1 NAND2X1_724 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf1), .B(_4145_), .Y(_4146_) );
OAI21X1 OAI21X1_1622 ( .gnd(gnd), .vdd(vdd), .A(_4146_), .B(_4144_), .C(raddr2_1_bF_buf9_), .Y(_4147_) );
OAI22X1 OAI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(_4140_), .B(_4141_), .C(_4147_), .D(_4143_), .Y(_4148_) );
AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_4148_), .B(_4033__bF_buf2), .C(_4132_), .D(_4138_), .Y(_4149_) );
OAI21X1 OAI21X1_1623 ( .gnd(gnd), .vdd(vdd), .A(_2530_), .B(raddr2_0_bF_buf22_), .C(raddr2_1_bF_buf8_), .Y(_4150_) );
AOI21X1 AOI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(regs_4__2_), .B(raddr2_0_bF_buf21_), .C(_4150_), .Y(_4151_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(regs_6__2_), .B(raddr2_0_bF_buf20_), .Y(_4152_) );
OAI21X1 OAI21X1_1624 ( .gnd(gnd), .vdd(vdd), .A(_2105_), .B(raddr2_0_bF_buf19_), .C(_4038__bF_buf0), .Y(_4153_) );
OAI21X1 OAI21X1_1625 ( .gnd(gnd), .vdd(vdd), .A(_4153_), .B(_4152_), .C(_4036__bF_buf0), .Y(_4154_) );
OAI21X1 OAI21X1_1626 ( .gnd(gnd), .vdd(vdd), .A(_2537_), .B(raddr2_0_bF_buf18_), .C(raddr2_1_bF_buf7_), .Y(_4155_) );
AOI21X1 AOI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(regs_0__2_), .B(raddr2_0_bF_buf17_), .C(_4155_), .Y(_4156_) );
NOR2X1 NOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf16_), .B(_2534_), .Y(_4157_) );
NAND2X1 NAND2X1_725 ( .gnd(gnd), .vdd(vdd), .A(regs_2__2_), .B(raddr2_0_bF_buf15_), .Y(_4158_) );
NAND2X1 NAND2X1_726 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf8), .B(_4158_), .Y(_4159_) );
OAI21X1 OAI21X1_1627 ( .gnd(gnd), .vdd(vdd), .A(_4159_), .B(_4157_), .C(raddr2_2_bF_buf10_), .Y(_4160_) );
OAI22X1 OAI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(_4156_), .B(_4160_), .C(_4154_), .D(_4151_), .Y(_4161_) );
NAND2X1 NAND2X1_727 ( .gnd(gnd), .vdd(vdd), .A(regs_10__2_), .B(raddr2_0_bF_buf14_), .Y(_4162_) );
OAI21X1 OAI21X1_1628 ( .gnd(gnd), .vdd(vdd), .A(_1906_), .B(raddr2_0_bF_buf13_), .C(_4162_), .Y(_4163_) );
NAND2X1 NAND2X1_728 ( .gnd(gnd), .vdd(vdd), .A(regs_8__2_), .B(raddr2_0_bF_buf12_), .Y(_4164_) );
OAI21X1 OAI21X1_1629 ( .gnd(gnd), .vdd(vdd), .A(_2004_), .B(raddr2_0_bF_buf11_), .C(_4164_), .Y(_4165_) );
MUX2X1 MUX2X1_321 ( .gnd(gnd), .vdd(vdd), .A(_4165_), .B(_4163_), .S(raddr2_1_bF_buf6_), .Y(_4166_) );
NAND2X1 NAND2X1_729 ( .gnd(gnd), .vdd(vdd), .A(regs_14__2_), .B(raddr2_0_bF_buf10_), .Y(_4167_) );
OAI21X1 OAI21X1_1630 ( .gnd(gnd), .vdd(vdd), .A(_1709_), .B(raddr2_0_bF_buf9_), .C(_4167_), .Y(_4168_) );
NAND2X1 NAND2X1_730 ( .gnd(gnd), .vdd(vdd), .A(regs_12__2_), .B(raddr2_0_bF_buf8_), .Y(_4169_) );
OAI21X1 OAI21X1_1631 ( .gnd(gnd), .vdd(vdd), .A(_1807_), .B(raddr2_0_bF_buf7_), .C(_4169_), .Y(_4170_) );
MUX2X1 MUX2X1_322 ( .gnd(gnd), .vdd(vdd), .A(_4170_), .B(_4168_), .S(raddr2_1_bF_buf5_), .Y(_4171_) );
MUX2X1 MUX2X1_323 ( .gnd(gnd), .vdd(vdd), .A(_4171_), .B(_4166_), .S(_4036__bF_buf8), .Y(_4172_) );
MUX2X1 MUX2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_4172_), .B(_4161_), .S(_4033__bF_buf1), .Y(_4173_) );
MUX2X1 MUX2X1_325 ( .gnd(gnd), .vdd(vdd), .A(_4173_), .B(_4149_), .S(raddr2_4_bF_buf2_), .Y(_5512__2_) );
NAND2X1 NAND2X1_731 ( .gnd(gnd), .vdd(vdd), .A(regs_22__3_), .B(raddr2_0_bF_buf6_), .Y(_4174_) );
OAI21X1 OAI21X1_1632 ( .gnd(gnd), .vdd(vdd), .A(_1316_), .B(raddr2_0_bF_buf5_), .C(_4174_), .Y(_4175_) );
NAND2X1 NAND2X1_732 ( .gnd(gnd), .vdd(vdd), .A(regs_20__3_), .B(raddr2_0_bF_buf4_), .Y(_4176_) );
OAI21X1 OAI21X1_1633 ( .gnd(gnd), .vdd(vdd), .A(_1414_), .B(raddr2_0_bF_buf3_), .C(_4176_), .Y(_4177_) );
MUX2X1 MUX2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_4177_), .B(_4175_), .S(raddr2_1_bF_buf4_), .Y(_4178_) );
NAND2X1 NAND2X1_733 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf7), .B(_4178_), .Y(_4179_) );
NAND2X1 NAND2X1_734 ( .gnd(gnd), .vdd(vdd), .A(regs_18__3_), .B(raddr2_0_bF_buf2_), .Y(_4180_) );
OAI21X1 OAI21X1_1634 ( .gnd(gnd), .vdd(vdd), .A(_1513_), .B(raddr2_0_bF_buf1_), .C(_4180_), .Y(_4181_) );
NAND2X1 NAND2X1_735 ( .gnd(gnd), .vdd(vdd), .A(regs_16__3_), .B(raddr2_0_bF_buf0_), .Y(_4182_) );
OAI21X1 OAI21X1_1635 ( .gnd(gnd), .vdd(vdd), .A(_1611_), .B(raddr2_0_bF_buf96_), .C(_4182_), .Y(_4183_) );
MUX2X1 MUX2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_4183_), .B(_4181_), .S(raddr2_1_bF_buf3_), .Y(_4184_) );
AOI21X1 AOI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(raddr2_2_bF_buf9_), .B(_4184_), .C(_4033__bF_buf0), .Y(_4185_) );
OAI21X1 OAI21X1_1636 ( .gnd(gnd), .vdd(vdd), .A(_1149_), .B(raddr2_0_bF_buf95_), .C(raddr2_2_bF_buf8_), .Y(_4186_) );
AOI21X1 AOI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(regs_26__3_), .B(raddr2_0_bF_buf94_), .C(_4186_), .Y(_4187_) );
OAI21X1 OAI21X1_1637 ( .gnd(gnd), .vdd(vdd), .A(regs_30__3_), .B(raddr2_2_bF_buf7_), .C(_4038__bF_buf7), .Y(_4188_) );
OAI21X1 OAI21X1_1638 ( .gnd(gnd), .vdd(vdd), .A(_2599_), .B(raddr2_0_bF_buf93_), .C(raddr2_2_bF_buf6_), .Y(_4189_) );
AOI21X1 AOI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(regs_24__3_), .B(raddr2_0_bF_buf92_), .C(_4189_), .Y(_4190_) );
NOR2X1 NOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf91_), .B(_2593_), .Y(_4191_) );
NAND2X1 NAND2X1_736 ( .gnd(gnd), .vdd(vdd), .A(regs_28__3_), .B(raddr2_0_bF_buf90_), .Y(_4192_) );
NAND2X1 NAND2X1_737 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf6), .B(_4192_), .Y(_4193_) );
OAI21X1 OAI21X1_1639 ( .gnd(gnd), .vdd(vdd), .A(_4193_), .B(_4191_), .C(raddr2_1_bF_buf2_), .Y(_4194_) );
OAI22X1 OAI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(_4187_), .B(_4188_), .C(_4194_), .D(_4190_), .Y(_4195_) );
AOI22X1 AOI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_4195_), .B(_4033__bF_buf7), .C(_4179_), .D(_4185_), .Y(_4196_) );
OAI21X1 OAI21X1_1640 ( .gnd(gnd), .vdd(vdd), .A(_2554_), .B(raddr2_0_bF_buf89_), .C(raddr2_1_bF_buf1_), .Y(_4197_) );
AOI21X1 AOI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(regs_4__3_), .B(raddr2_0_bF_buf88_), .C(_4197_), .Y(_4198_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(regs_6__3_), .B(raddr2_0_bF_buf87_), .Y(_4199_) );
OAI21X1 OAI21X1_1641 ( .gnd(gnd), .vdd(vdd), .A(_2107_), .B(raddr2_0_bF_buf86_), .C(_4038__bF_buf6), .Y(_4200_) );
OAI21X1 OAI21X1_1642 ( .gnd(gnd), .vdd(vdd), .A(_4200_), .B(_4199_), .C(_4036__bF_buf5), .Y(_4201_) );
OAI21X1 OAI21X1_1643 ( .gnd(gnd), .vdd(vdd), .A(_2560_), .B(raddr2_0_bF_buf85_), .C(raddr2_1_bF_buf0_), .Y(_4202_) );
AOI21X1 AOI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(regs_0__3_), .B(raddr2_0_bF_buf84_), .C(_4202_), .Y(_4203_) );
NOR2X1 NOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf83_), .B(_2563_), .Y(_4204_) );
NAND2X1 NAND2X1_738 ( .gnd(gnd), .vdd(vdd), .A(regs_2__3_), .B(raddr2_0_bF_buf82_), .Y(_4205_) );
NAND2X1 NAND2X1_739 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf5), .B(_4205_), .Y(_4206_) );
OAI21X1 OAI21X1_1644 ( .gnd(gnd), .vdd(vdd), .A(_4206_), .B(_4204_), .C(raddr2_2_bF_buf5_), .Y(_4207_) );
OAI22X1 OAI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(_4203_), .B(_4207_), .C(_4201_), .D(_4198_), .Y(_4208_) );
NAND2X1 NAND2X1_740 ( .gnd(gnd), .vdd(vdd), .A(regs_10__3_), .B(raddr2_0_bF_buf81_), .Y(_4209_) );
OAI21X1 OAI21X1_1645 ( .gnd(gnd), .vdd(vdd), .A(_1908_), .B(raddr2_0_bF_buf80_), .C(_4209_), .Y(_4210_) );
NAND2X1 NAND2X1_741 ( .gnd(gnd), .vdd(vdd), .A(regs_8__3_), .B(raddr2_0_bF_buf79_), .Y(_4211_) );
OAI21X1 OAI21X1_1646 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .B(raddr2_0_bF_buf78_), .C(_4211_), .Y(_4212_) );
MUX2X1 MUX2X1_328 ( .gnd(gnd), .vdd(vdd), .A(_4212_), .B(_4210_), .S(raddr2_1_bF_buf14_bF_buf1_), .Y(_4213_) );
NAND2X1 NAND2X1_742 ( .gnd(gnd), .vdd(vdd), .A(regs_14__3_), .B(raddr2_0_bF_buf77_), .Y(_4214_) );
OAI21X1 OAI21X1_1647 ( .gnd(gnd), .vdd(vdd), .A(_1711_), .B(raddr2_0_bF_buf76_), .C(_4214_), .Y(_4215_) );
NAND2X1 NAND2X1_743 ( .gnd(gnd), .vdd(vdd), .A(regs_12__3_), .B(raddr2_0_bF_buf75_), .Y(_4216_) );
OAI21X1 OAI21X1_1648 ( .gnd(gnd), .vdd(vdd), .A(_1809_), .B(raddr2_0_bF_buf74_), .C(_4216_), .Y(_4217_) );
MUX2X1 MUX2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_4217_), .B(_4215_), .S(raddr2_1_bF_buf13_bF_buf1_), .Y(_4218_) );
MUX2X1 MUX2X1_330 ( .gnd(gnd), .vdd(vdd), .A(_4218_), .B(_4213_), .S(_4036__bF_buf4), .Y(_4219_) );
MUX2X1 MUX2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_4219_), .B(_4208_), .S(_4033__bF_buf6), .Y(_4220_) );
MUX2X1 MUX2X1_332 ( .gnd(gnd), .vdd(vdd), .A(_4220_), .B(_4196_), .S(raddr2_4_bF_buf1_), .Y(_5512__3_) );
OAI21X1 OAI21X1_1649 ( .gnd(gnd), .vdd(vdd), .A(_2605_), .B(raddr2_0_bF_buf73_), .C(raddr2_1_bF_buf12_bF_buf1_), .Y(_4221_) );
AOI21X1 AOI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(regs_4__4_), .B(raddr2_0_bF_buf72_), .C(_4221_), .Y(_4222_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(regs_6__4_), .B(raddr2_0_bF_buf71_), .Y(_4223_) );
OAI21X1 OAI21X1_1650 ( .gnd(gnd), .vdd(vdd), .A(_2109_), .B(raddr2_0_bF_buf70_), .C(_4038__bF_buf4), .Y(_4224_) );
OAI21X1 OAI21X1_1651 ( .gnd(gnd), .vdd(vdd), .A(_4224_), .B(_4223_), .C(_4036__bF_buf3), .Y(_4225_) );
OAI21X1 OAI21X1_1652 ( .gnd(gnd), .vdd(vdd), .A(_2611_), .B(raddr2_0_bF_buf69_), .C(raddr2_1_bF_buf11_), .Y(_4226_) );
AOI21X1 AOI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(regs_0__4_), .B(raddr2_0_bF_buf68_), .C(_4226_), .Y(_4227_) );
NOR2X1 NOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf67_), .B(_2614_), .Y(_4228_) );
NAND2X1 NAND2X1_744 ( .gnd(gnd), .vdd(vdd), .A(regs_2__4_), .B(raddr2_0_bF_buf66_), .Y(_4229_) );
NAND2X1 NAND2X1_745 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf3), .B(_4229_), .Y(_4230_) );
OAI21X1 OAI21X1_1653 ( .gnd(gnd), .vdd(vdd), .A(_4230_), .B(_4228_), .C(raddr2_2_bF_buf4_), .Y(_4231_) );
OAI22X1 OAI22X1_61 ( .gnd(gnd), .vdd(vdd), .A(_4227_), .B(_4231_), .C(_4225_), .D(_4222_), .Y(_4232_) );
NAND2X1 NAND2X1_746 ( .gnd(gnd), .vdd(vdd), .A(regs_10__4_), .B(raddr2_0_bF_buf65_), .Y(_4233_) );
OAI21X1 OAI21X1_1654 ( .gnd(gnd), .vdd(vdd), .A(_1910_), .B(raddr2_0_bF_buf64_), .C(_4233_), .Y(_4234_) );
NAND2X1 NAND2X1_747 ( .gnd(gnd), .vdd(vdd), .A(regs_8__4_), .B(raddr2_0_bF_buf63_), .Y(_4235_) );
OAI21X1 OAI21X1_1655 ( .gnd(gnd), .vdd(vdd), .A(_2008_), .B(raddr2_0_bF_buf62_), .C(_4235_), .Y(_4236_) );
MUX2X1 MUX2X1_333 ( .gnd(gnd), .vdd(vdd), .A(_4236_), .B(_4234_), .S(raddr2_1_bF_buf10_), .Y(_4237_) );
NAND2X1 NAND2X1_748 ( .gnd(gnd), .vdd(vdd), .A(regs_14__4_), .B(raddr2_0_bF_buf61_), .Y(_4238_) );
OAI21X1 OAI21X1_1656 ( .gnd(gnd), .vdd(vdd), .A(_1713_), .B(raddr2_0_bF_buf60_), .C(_4238_), .Y(_4239_) );
NAND2X1 NAND2X1_749 ( .gnd(gnd), .vdd(vdd), .A(regs_12__4_), .B(raddr2_0_bF_buf59_), .Y(_4240_) );
OAI21X1 OAI21X1_1657 ( .gnd(gnd), .vdd(vdd), .A(_1811_), .B(raddr2_0_bF_buf58_), .C(_4240_), .Y(_4241_) );
MUX2X1 MUX2X1_334 ( .gnd(gnd), .vdd(vdd), .A(_4241_), .B(_4239_), .S(raddr2_1_bF_buf9_), .Y(_4242_) );
MUX2X1 MUX2X1_335 ( .gnd(gnd), .vdd(vdd), .A(_4242_), .B(_4237_), .S(_4036__bF_buf2), .Y(_4243_) );
MUX2X1 MUX2X1_336 ( .gnd(gnd), .vdd(vdd), .A(_4243_), .B(_4232_), .S(_4033__bF_buf5), .Y(_4244_) );
OAI21X1 OAI21X1_1658 ( .gnd(gnd), .vdd(vdd), .A(_1613_), .B(raddr2_0_bF_buf57_), .C(raddr2_1_bF_buf8_), .Y(_4245_) );
AOI21X1 AOI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(regs_16__4_), .B(raddr2_0_bF_buf56_), .C(_4245_), .Y(_4246_) );
NOR2X1 NOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf55_), .B(_1515_), .Y(_4247_) );
NAND2X1 NAND2X1_750 ( .gnd(gnd), .vdd(vdd), .A(regs_18__4_), .B(raddr2_0_bF_buf54_), .Y(_4248_) );
NAND2X1 NAND2X1_751 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf2), .B(_4248_), .Y(_4249_) );
OAI21X1 OAI21X1_1659 ( .gnd(gnd), .vdd(vdd), .A(_4249_), .B(_4247_), .C(raddr2_2_bF_buf3_), .Y(_4250_) );
OAI21X1 OAI21X1_1660 ( .gnd(gnd), .vdd(vdd), .A(_1416_), .B(raddr2_0_bF_buf53_), .C(raddr2_1_bF_buf7_), .Y(_4251_) );
AOI21X1 AOI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(regs_20__4_), .B(raddr2_0_bF_buf52_), .C(_4251_), .Y(_4252_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(regs_22__4_), .B(raddr2_0_bF_buf51_), .Y(_4253_) );
OAI21X1 OAI21X1_1661 ( .gnd(gnd), .vdd(vdd), .A(_1318_), .B(raddr2_0_bF_buf50_), .C(_4038__bF_buf1), .Y(_4254_) );
OAI21X1 OAI21X1_1662 ( .gnd(gnd), .vdd(vdd), .A(_4254_), .B(_4253_), .C(_4036__bF_buf1), .Y(_4255_) );
OAI22X1 OAI22X1_62 ( .gnd(gnd), .vdd(vdd), .A(_4246_), .B(_4250_), .C(_4255_), .D(_4252_), .Y(_4256_) );
NAND2X1 NAND2X1_752 ( .gnd(gnd), .vdd(vdd), .A(regs_28__4_), .B(raddr2_0_bF_buf49_), .Y(_4257_) );
OAI21X1 OAI21X1_1663 ( .gnd(gnd), .vdd(vdd), .A(_2644_), .B(raddr2_0_bF_buf48_), .C(_4257_), .Y(_4258_) );
MUX2X1 MUX2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_4258_), .B(regs_30__4_), .S(raddr2_1_bF_buf6_), .Y(_4259_) );
NAND2X1 NAND2X1_753 ( .gnd(gnd), .vdd(vdd), .A(regs_26__4_), .B(raddr2_0_bF_buf47_), .Y(_4260_) );
OAI21X1 OAI21X1_1664 ( .gnd(gnd), .vdd(vdd), .A(_1151_), .B(raddr2_0_bF_buf46_), .C(_4260_), .Y(_4261_) );
NAND2X1 NAND2X1_754 ( .gnd(gnd), .vdd(vdd), .A(regs_24__4_), .B(raddr2_0_bF_buf45_), .Y(_4262_) );
OAI21X1 OAI21X1_1665 ( .gnd(gnd), .vdd(vdd), .A(_2650_), .B(raddr2_0_bF_buf44_), .C(_4262_), .Y(_4263_) );
MUX2X1 MUX2X1_338 ( .gnd(gnd), .vdd(vdd), .A(_4263_), .B(_4261_), .S(raddr2_1_bF_buf5_), .Y(_4264_) );
MUX2X1 MUX2X1_339 ( .gnd(gnd), .vdd(vdd), .A(_4264_), .B(_4259_), .S(raddr2_2_bF_buf2_), .Y(_4265_) );
MUX2X1 MUX2X1_340 ( .gnd(gnd), .vdd(vdd), .A(_4265_), .B(_4256_), .S(_4033__bF_buf4), .Y(_4266_) );
MUX2X1 MUX2X1_341 ( .gnd(gnd), .vdd(vdd), .A(_4244_), .B(_4266_), .S(raddr2_4_bF_buf0_), .Y(_5512__4_) );
OAI21X1 OAI21X1_1666 ( .gnd(gnd), .vdd(vdd), .A(_1418_), .B(raddr2_0_bF_buf43_), .C(raddr2_1_bF_buf4_), .Y(_4267_) );
AOI21X1 AOI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(regs_20__5_), .B(raddr2_0_bF_buf42_), .C(_4267_), .Y(_4268_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(regs_22__5_), .B(raddr2_0_bF_buf41_), .Y(_4269_) );
OAI21X1 OAI21X1_1667 ( .gnd(gnd), .vdd(vdd), .A(_1320_), .B(raddr2_0_bF_buf40_), .C(_4038__bF_buf0), .Y(_4270_) );
OAI21X1 OAI21X1_1668 ( .gnd(gnd), .vdd(vdd), .A(_4270_), .B(_4269_), .C(_4036__bF_buf0), .Y(_4271_) );
OAI21X1 OAI21X1_1669 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(raddr2_0_bF_buf39_), .C(raddr2_1_bF_buf3_), .Y(_4272_) );
AOI21X1 AOI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(regs_16__5_), .B(raddr2_0_bF_buf38_), .C(_4272_), .Y(_4273_) );
NOR2X1 NOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf37_), .B(_1517_), .Y(_4274_) );
NAND2X1 NAND2X1_755 ( .gnd(gnd), .vdd(vdd), .A(regs_18__5_), .B(raddr2_0_bF_buf36_), .Y(_4275_) );
NAND2X1 NAND2X1_756 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf8), .B(_4275_), .Y(_4276_) );
OAI21X1 OAI21X1_1670 ( .gnd(gnd), .vdd(vdd), .A(_4276_), .B(_4274_), .C(raddr2_2_bF_buf1_), .Y(_4277_) );
OAI22X1 OAI22X1_63 ( .gnd(gnd), .vdd(vdd), .A(_4273_), .B(_4277_), .C(_4271_), .D(_4268_), .Y(_4278_) );
NAND2X1 NAND2X1_757 ( .gnd(gnd), .vdd(vdd), .A(regs_28__5_), .B(raddr2_0_bF_buf35_), .Y(_4279_) );
OAI21X1 OAI21X1_1671 ( .gnd(gnd), .vdd(vdd), .A(_2668_), .B(raddr2_0_bF_buf34_), .C(_4279_), .Y(_4280_) );
MUX2X1 MUX2X1_342 ( .gnd(gnd), .vdd(vdd), .A(_4280_), .B(regs_30__5_), .S(raddr2_1_bF_buf2_), .Y(_4281_) );
NAND2X1 NAND2X1_758 ( .gnd(gnd), .vdd(vdd), .A(regs_26__5_), .B(raddr2_0_bF_buf33_), .Y(_4282_) );
OAI21X1 OAI21X1_1672 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(raddr2_0_bF_buf32_), .C(_4282_), .Y(_4283_) );
NAND2X1 NAND2X1_759 ( .gnd(gnd), .vdd(vdd), .A(regs_24__5_), .B(raddr2_0_bF_buf31_), .Y(_4284_) );
OAI21X1 OAI21X1_1673 ( .gnd(gnd), .vdd(vdd), .A(_2674_), .B(raddr2_0_bF_buf30_), .C(_4284_), .Y(_4285_) );
MUX2X1 MUX2X1_343 ( .gnd(gnd), .vdd(vdd), .A(_4285_), .B(_4283_), .S(raddr2_1_bF_buf1_), .Y(_4286_) );
MUX2X1 MUX2X1_344 ( .gnd(gnd), .vdd(vdd), .A(_4286_), .B(_4281_), .S(raddr2_2_bF_buf0_), .Y(_4287_) );
MUX2X1 MUX2X1_345 ( .gnd(gnd), .vdd(vdd), .A(_4287_), .B(_4278_), .S(_4033__bF_buf3), .Y(_4288_) );
NAND2X1 NAND2X1_760 ( .gnd(gnd), .vdd(vdd), .A(regs_6__5_), .B(raddr2_0_bF_buf29_), .Y(_4289_) );
OAI21X1 OAI21X1_1674 ( .gnd(gnd), .vdd(vdd), .A(_2111_), .B(raddr2_0_bF_buf28_), .C(_4289_), .Y(_4290_) );
NAND2X1 NAND2X1_761 ( .gnd(gnd), .vdd(vdd), .A(regs_4__5_), .B(raddr2_0_bF_buf27_), .Y(_4291_) );
OAI21X1 OAI21X1_1675 ( .gnd(gnd), .vdd(vdd), .A(_2682_), .B(raddr2_0_bF_buf26_), .C(_4291_), .Y(_4292_) );
MUX2X1 MUX2X1_346 ( .gnd(gnd), .vdd(vdd), .A(_4292_), .B(_4290_), .S(raddr2_1_bF_buf0_), .Y(_4293_) );
NAND2X1 NAND2X1_762 ( .gnd(gnd), .vdd(vdd), .A(regs_2__5_), .B(raddr2_0_bF_buf25_), .Y(_4294_) );
OAI21X1 OAI21X1_1676 ( .gnd(gnd), .vdd(vdd), .A(_2686_), .B(raddr2_0_bF_buf24_), .C(_4294_), .Y(_4295_) );
NAND2X1 NAND2X1_763 ( .gnd(gnd), .vdd(vdd), .A(regs_0__5_), .B(raddr2_0_bF_buf23_), .Y(_4296_) );
OAI21X1 OAI21X1_1677 ( .gnd(gnd), .vdd(vdd), .A(_2689_), .B(raddr2_0_bF_buf22_), .C(_4296_), .Y(_4297_) );
MUX2X1 MUX2X1_347 ( .gnd(gnd), .vdd(vdd), .A(_4297_), .B(_4295_), .S(raddr2_1_bF_buf14_bF_buf0_), .Y(_4298_) );
MUX2X1 MUX2X1_348 ( .gnd(gnd), .vdd(vdd), .A(_4298_), .B(_4293_), .S(raddr2_2_bF_buf10_), .Y(_4299_) );
NAND2X1 NAND2X1_764 ( .gnd(gnd), .vdd(vdd), .A(regs_14__5_), .B(raddr2_0_bF_buf21_), .Y(_4300_) );
OAI21X1 OAI21X1_1678 ( .gnd(gnd), .vdd(vdd), .A(_1715_), .B(raddr2_0_bF_buf20_), .C(_4300_), .Y(_4301_) );
NAND2X1 NAND2X1_765 ( .gnd(gnd), .vdd(vdd), .A(regs_12__5_), .B(raddr2_0_bF_buf19_), .Y(_4302_) );
OAI21X1 OAI21X1_1679 ( .gnd(gnd), .vdd(vdd), .A(_1813_), .B(raddr2_0_bF_buf18_), .C(_4302_), .Y(_4303_) );
MUX2X1 MUX2X1_349 ( .gnd(gnd), .vdd(vdd), .A(_4303_), .B(_4301_), .S(raddr2_1_bF_buf13_bF_buf0_), .Y(_4304_) );
NAND2X1 NAND2X1_766 ( .gnd(gnd), .vdd(vdd), .A(regs_10__5_), .B(raddr2_0_bF_buf17_), .Y(_4305_) );
OAI21X1 OAI21X1_1680 ( .gnd(gnd), .vdd(vdd), .A(_1912_), .B(raddr2_0_bF_buf16_), .C(_4305_), .Y(_4306_) );
NAND2X1 NAND2X1_767 ( .gnd(gnd), .vdd(vdd), .A(regs_8__5_), .B(raddr2_0_bF_buf15_), .Y(_4307_) );
OAI21X1 OAI21X1_1681 ( .gnd(gnd), .vdd(vdd), .A(_2010_), .B(raddr2_0_bF_buf14_), .C(_4307_), .Y(_4308_) );
MUX2X1 MUX2X1_350 ( .gnd(gnd), .vdd(vdd), .A(_4308_), .B(_4306_), .S(raddr2_1_bF_buf12_bF_buf0_), .Y(_4309_) );
MUX2X1 MUX2X1_351 ( .gnd(gnd), .vdd(vdd), .A(_4309_), .B(_4304_), .S(raddr2_2_bF_buf9_), .Y(_4310_) );
MUX2X1 MUX2X1_352 ( .gnd(gnd), .vdd(vdd), .A(_4310_), .B(_4299_), .S(_4033__bF_buf2), .Y(_4311_) );
MUX2X1 MUX2X1_353 ( .gnd(gnd), .vdd(vdd), .A(_4311_), .B(_4288_), .S(raddr2_4_bF_buf4_), .Y(_5512__5_) );
OAI21X1 OAI21X1_1682 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(raddr2_0_bF_buf13_), .C(raddr2_1_bF_buf11_), .Y(_4312_) );
AOI21X1 AOI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(regs_20__6_), .B(raddr2_0_bF_buf12_), .C(_4312_), .Y(_4313_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(regs_22__6_), .B(raddr2_0_bF_buf11_), .Y(_4314_) );
OAI21X1 OAI21X1_1683 ( .gnd(gnd), .vdd(vdd), .A(_1322_), .B(raddr2_0_bF_buf10_), .C(_4038__bF_buf7), .Y(_4315_) );
OAI21X1 OAI21X1_1684 ( .gnd(gnd), .vdd(vdd), .A(_4315_), .B(_4314_), .C(_4036__bF_buf8), .Y(_4316_) );
OAI21X1 OAI21X1_1685 ( .gnd(gnd), .vdd(vdd), .A(_1617_), .B(raddr2_0_bF_buf9_), .C(raddr2_1_bF_buf10_), .Y(_4317_) );
AOI21X1 AOI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(regs_16__6_), .B(raddr2_0_bF_buf8_), .C(_4317_), .Y(_4318_) );
NOR2X1 NOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf7_), .B(_1519_), .Y(_4319_) );
NAND2X1 NAND2X1_768 ( .gnd(gnd), .vdd(vdd), .A(regs_18__6_), .B(raddr2_0_bF_buf6_), .Y(_4320_) );
NAND2X1 NAND2X1_769 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf6), .B(_4320_), .Y(_4321_) );
OAI21X1 OAI21X1_1686 ( .gnd(gnd), .vdd(vdd), .A(_4321_), .B(_4319_), .C(raddr2_2_bF_buf8_), .Y(_4322_) );
OAI22X1 OAI22X1_64 ( .gnd(gnd), .vdd(vdd), .A(_4318_), .B(_4322_), .C(_4316_), .D(_4313_), .Y(_4323_) );
NAND2X1 NAND2X1_770 ( .gnd(gnd), .vdd(vdd), .A(regs_28__6_), .B(raddr2_0_bF_buf5_), .Y(_4324_) );
OAI21X1 OAI21X1_1687 ( .gnd(gnd), .vdd(vdd), .A(_2718_), .B(raddr2_0_bF_buf4_), .C(_4324_), .Y(_4325_) );
MUX2X1 MUX2X1_354 ( .gnd(gnd), .vdd(vdd), .A(_4325_), .B(regs_30__6_), .S(raddr2_1_bF_buf9_), .Y(_4326_) );
NAND2X1 NAND2X1_771 ( .gnd(gnd), .vdd(vdd), .A(regs_26__6_), .B(raddr2_0_bF_buf3_), .Y(_4327_) );
OAI21X1 OAI21X1_1688 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .B(raddr2_0_bF_buf2_), .C(_4327_), .Y(_4328_) );
NAND2X1 NAND2X1_772 ( .gnd(gnd), .vdd(vdd), .A(regs_24__6_), .B(raddr2_0_bF_buf1_), .Y(_4329_) );
OAI21X1 OAI21X1_1689 ( .gnd(gnd), .vdd(vdd), .A(_2724_), .B(raddr2_0_bF_buf0_), .C(_4329_), .Y(_4330_) );
MUX2X1 MUX2X1_355 ( .gnd(gnd), .vdd(vdd), .A(_4330_), .B(_4328_), .S(raddr2_1_bF_buf8_), .Y(_4331_) );
MUX2X1 MUX2X1_356 ( .gnd(gnd), .vdd(vdd), .A(_4331_), .B(_4326_), .S(raddr2_2_bF_buf7_), .Y(_4332_) );
MUX2X1 MUX2X1_357 ( .gnd(gnd), .vdd(vdd), .A(_4332_), .B(_4323_), .S(_4033__bF_buf1), .Y(_4333_) );
NAND2X1 NAND2X1_773 ( .gnd(gnd), .vdd(vdd), .A(regs_6__6_), .B(raddr2_0_bF_buf96_), .Y(_4334_) );
OAI21X1 OAI21X1_1690 ( .gnd(gnd), .vdd(vdd), .A(_2113_), .B(raddr2_0_bF_buf95_), .C(_4334_), .Y(_4335_) );
NAND2X1 NAND2X1_774 ( .gnd(gnd), .vdd(vdd), .A(regs_4__6_), .B(raddr2_0_bF_buf94_), .Y(_4336_) );
OAI21X1 OAI21X1_1691 ( .gnd(gnd), .vdd(vdd), .A(_2732_), .B(raddr2_0_bF_buf93_), .C(_4336_), .Y(_4337_) );
MUX2X1 MUX2X1_358 ( .gnd(gnd), .vdd(vdd), .A(_4337_), .B(_4335_), .S(raddr2_1_bF_buf7_), .Y(_4338_) );
NAND2X1 NAND2X1_775 ( .gnd(gnd), .vdd(vdd), .A(regs_2__6_), .B(raddr2_0_bF_buf92_), .Y(_4339_) );
OAI21X1 OAI21X1_1692 ( .gnd(gnd), .vdd(vdd), .A(_2736_), .B(raddr2_0_bF_buf91_), .C(_4339_), .Y(_4340_) );
NAND2X1 NAND2X1_776 ( .gnd(gnd), .vdd(vdd), .A(regs_0__6_), .B(raddr2_0_bF_buf90_), .Y(_4341_) );
OAI21X1 OAI21X1_1693 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(raddr2_0_bF_buf89_), .C(_4341_), .Y(_4342_) );
MUX2X1 MUX2X1_359 ( .gnd(gnd), .vdd(vdd), .A(_4342_), .B(_4340_), .S(raddr2_1_bF_buf6_), .Y(_4343_) );
MUX2X1 MUX2X1_360 ( .gnd(gnd), .vdd(vdd), .A(_4343_), .B(_4338_), .S(raddr2_2_bF_buf6_), .Y(_4344_) );
NAND2X1 NAND2X1_777 ( .gnd(gnd), .vdd(vdd), .A(regs_14__6_), .B(raddr2_0_bF_buf88_), .Y(_4345_) );
OAI21X1 OAI21X1_1694 ( .gnd(gnd), .vdd(vdd), .A(_1717_), .B(raddr2_0_bF_buf87_), .C(_4345_), .Y(_4346_) );
NAND2X1 NAND2X1_778 ( .gnd(gnd), .vdd(vdd), .A(regs_12__6_), .B(raddr2_0_bF_buf86_), .Y(_4347_) );
OAI21X1 OAI21X1_1695 ( .gnd(gnd), .vdd(vdd), .A(_1815_), .B(raddr2_0_bF_buf85_), .C(_4347_), .Y(_4348_) );
MUX2X1 MUX2X1_361 ( .gnd(gnd), .vdd(vdd), .A(_4348_), .B(_4346_), .S(raddr2_1_bF_buf5_), .Y(_4349_) );
NAND2X1 NAND2X1_779 ( .gnd(gnd), .vdd(vdd), .A(regs_10__6_), .B(raddr2_0_bF_buf84_), .Y(_4350_) );
OAI21X1 OAI21X1_1696 ( .gnd(gnd), .vdd(vdd), .A(_1914_), .B(raddr2_0_bF_buf83_), .C(_4350_), .Y(_4351_) );
NAND2X1 NAND2X1_780 ( .gnd(gnd), .vdd(vdd), .A(regs_8__6_), .B(raddr2_0_bF_buf82_), .Y(_4352_) );
OAI21X1 OAI21X1_1697 ( .gnd(gnd), .vdd(vdd), .A(_2012_), .B(raddr2_0_bF_buf81_), .C(_4352_), .Y(_4353_) );
MUX2X1 MUX2X1_362 ( .gnd(gnd), .vdd(vdd), .A(_4353_), .B(_4351_), .S(raddr2_1_bF_buf4_), .Y(_4354_) );
MUX2X1 MUX2X1_363 ( .gnd(gnd), .vdd(vdd), .A(_4354_), .B(_4349_), .S(raddr2_2_bF_buf5_), .Y(_4355_) );
MUX2X1 MUX2X1_364 ( .gnd(gnd), .vdd(vdd), .A(_4355_), .B(_4344_), .S(_4033__bF_buf0), .Y(_4356_) );
MUX2X1 MUX2X1_365 ( .gnd(gnd), .vdd(vdd), .A(_4356_), .B(_4333_), .S(raddr2_4_bF_buf3_), .Y(_5512__6_) );
NAND2X1 NAND2X1_781 ( .gnd(gnd), .vdd(vdd), .A(regs_22__7_), .B(raddr2_0_bF_buf80_), .Y(_4357_) );
OAI21X1 OAI21X1_1698 ( .gnd(gnd), .vdd(vdd), .A(_1324_), .B(raddr2_0_bF_buf79_), .C(_4357_), .Y(_4358_) );
NAND2X1 NAND2X1_782 ( .gnd(gnd), .vdd(vdd), .A(regs_20__7_), .B(raddr2_0_bF_buf78_), .Y(_4359_) );
OAI21X1 OAI21X1_1699 ( .gnd(gnd), .vdd(vdd), .A(_1422_), .B(raddr2_0_bF_buf77_), .C(_4359_), .Y(_4360_) );
MUX2X1 MUX2X1_366 ( .gnd(gnd), .vdd(vdd), .A(_4360_), .B(_4358_), .S(raddr2_1_bF_buf3_), .Y(_4361_) );
NAND2X1 NAND2X1_783 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf7), .B(_4361_), .Y(_4362_) );
NAND2X1 NAND2X1_784 ( .gnd(gnd), .vdd(vdd), .A(regs_18__7_), .B(raddr2_0_bF_buf76_), .Y(_4363_) );
OAI21X1 OAI21X1_1700 ( .gnd(gnd), .vdd(vdd), .A(_1521_), .B(raddr2_0_bF_buf75_), .C(_4363_), .Y(_4364_) );
NAND2X1 NAND2X1_785 ( .gnd(gnd), .vdd(vdd), .A(regs_16__7_), .B(raddr2_0_bF_buf74_), .Y(_4365_) );
OAI21X1 OAI21X1_1701 ( .gnd(gnd), .vdd(vdd), .A(_1619_), .B(raddr2_0_bF_buf73_), .C(_4365_), .Y(_4366_) );
MUX2X1 MUX2X1_367 ( .gnd(gnd), .vdd(vdd), .A(_4366_), .B(_4364_), .S(raddr2_1_bF_buf2_), .Y(_4367_) );
AOI21X1 AOI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(raddr2_2_bF_buf4_), .B(_4367_), .C(_4033__bF_buf7), .Y(_4368_) );
OAI21X1 OAI21X1_1702 ( .gnd(gnd), .vdd(vdd), .A(_1157_), .B(raddr2_0_bF_buf72_), .C(raddr2_2_bF_buf3_), .Y(_4369_) );
AOI21X1 AOI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(regs_26__7_), .B(raddr2_0_bF_buf71_), .C(_4369_), .Y(_4370_) );
OAI21X1 OAI21X1_1703 ( .gnd(gnd), .vdd(vdd), .A(regs_30__7_), .B(raddr2_2_bF_buf2_), .C(_4038__bF_buf5), .Y(_4371_) );
OAI21X1 OAI21X1_1704 ( .gnd(gnd), .vdd(vdd), .A(_2771_), .B(raddr2_0_bF_buf70_), .C(raddr2_2_bF_buf1_), .Y(_4372_) );
AOI21X1 AOI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(regs_24__7_), .B(raddr2_0_bF_buf69_), .C(_4372_), .Y(_4373_) );
NOR2X1 NOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf68_), .B(_2774_), .Y(_4374_) );
NAND2X1 NAND2X1_786 ( .gnd(gnd), .vdd(vdd), .A(regs_28__7_), .B(raddr2_0_bF_buf67_), .Y(_4375_) );
NAND2X1 NAND2X1_787 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf6), .B(_4375_), .Y(_4376_) );
OAI21X1 OAI21X1_1705 ( .gnd(gnd), .vdd(vdd), .A(_4376_), .B(_4374_), .C(raddr2_1_bF_buf1_), .Y(_4377_) );
OAI22X1 OAI22X1_65 ( .gnd(gnd), .vdd(vdd), .A(_4370_), .B(_4371_), .C(_4377_), .D(_4373_), .Y(_4378_) );
AOI22X1 AOI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_4378_), .B(_4033__bF_buf6), .C(_4362_), .D(_4368_), .Y(_4379_) );
OAI21X1 OAI21X1_1706 ( .gnd(gnd), .vdd(vdd), .A(_2781_), .B(raddr2_0_bF_buf66_), .C(raddr2_1_bF_buf0_), .Y(_4380_) );
AOI21X1 AOI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(regs_4__7_), .B(raddr2_0_bF_buf65_), .C(_4380_), .Y(_4381_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(regs_6__7_), .B(raddr2_0_bF_buf64_), .Y(_4382_) );
OAI21X1 OAI21X1_1707 ( .gnd(gnd), .vdd(vdd), .A(_2115_), .B(raddr2_0_bF_buf63_), .C(_4038__bF_buf4), .Y(_4383_) );
OAI21X1 OAI21X1_1708 ( .gnd(gnd), .vdd(vdd), .A(_4383_), .B(_4382_), .C(_4036__bF_buf5), .Y(_4384_) );
OAI21X1 OAI21X1_1709 ( .gnd(gnd), .vdd(vdd), .A(_2787_), .B(raddr2_0_bF_buf62_), .C(raddr2_1_bF_buf14_bF_buf3_), .Y(_4385_) );
AOI21X1 AOI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(regs_0__7_), .B(raddr2_0_bF_buf61_), .C(_4385_), .Y(_4386_) );
NOR2X1 NOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf60_), .B(_2790_), .Y(_4387_) );
NAND2X1 NAND2X1_788 ( .gnd(gnd), .vdd(vdd), .A(regs_2__7_), .B(raddr2_0_bF_buf59_), .Y(_4388_) );
NAND2X1 NAND2X1_789 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf3), .B(_4388_), .Y(_4389_) );
OAI21X1 OAI21X1_1710 ( .gnd(gnd), .vdd(vdd), .A(_4389_), .B(_4387_), .C(raddr2_2_bF_buf0_), .Y(_4390_) );
OAI22X1 OAI22X1_66 ( .gnd(gnd), .vdd(vdd), .A(_4386_), .B(_4390_), .C(_4384_), .D(_4381_), .Y(_4391_) );
NAND2X1 NAND2X1_790 ( .gnd(gnd), .vdd(vdd), .A(regs_10__7_), .B(raddr2_0_bF_buf58_), .Y(_4392_) );
OAI21X1 OAI21X1_1711 ( .gnd(gnd), .vdd(vdd), .A(_1916_), .B(raddr2_0_bF_buf57_), .C(_4392_), .Y(_4393_) );
NAND2X1 NAND2X1_791 ( .gnd(gnd), .vdd(vdd), .A(regs_8__7_), .B(raddr2_0_bF_buf56_), .Y(_4394_) );
OAI21X1 OAI21X1_1712 ( .gnd(gnd), .vdd(vdd), .A(_2014_), .B(raddr2_0_bF_buf55_), .C(_4394_), .Y(_4395_) );
MUX2X1 MUX2X1_368 ( .gnd(gnd), .vdd(vdd), .A(_4395_), .B(_4393_), .S(raddr2_1_bF_buf13_bF_buf3_), .Y(_4396_) );
NAND2X1 NAND2X1_792 ( .gnd(gnd), .vdd(vdd), .A(regs_14__7_), .B(raddr2_0_bF_buf54_), .Y(_4397_) );
OAI21X1 OAI21X1_1713 ( .gnd(gnd), .vdd(vdd), .A(_1719_), .B(raddr2_0_bF_buf53_), .C(_4397_), .Y(_4398_) );
NAND2X1 NAND2X1_793 ( .gnd(gnd), .vdd(vdd), .A(regs_12__7_), .B(raddr2_0_bF_buf52_), .Y(_4399_) );
OAI21X1 OAI21X1_1714 ( .gnd(gnd), .vdd(vdd), .A(_1817_), .B(raddr2_0_bF_buf51_), .C(_4399_), .Y(_4400_) );
MUX2X1 MUX2X1_369 ( .gnd(gnd), .vdd(vdd), .A(_4400_), .B(_4398_), .S(raddr2_1_bF_buf12_bF_buf3_), .Y(_4401_) );
MUX2X1 MUX2X1_370 ( .gnd(gnd), .vdd(vdd), .A(_4401_), .B(_4396_), .S(_4036__bF_buf4), .Y(_4402_) );
MUX2X1 MUX2X1_371 ( .gnd(gnd), .vdd(vdd), .A(_4402_), .B(_4391_), .S(_4033__bF_buf5), .Y(_4403_) );
MUX2X1 MUX2X1_372 ( .gnd(gnd), .vdd(vdd), .A(_4403_), .B(_4379_), .S(raddr2_4_bF_buf2_), .Y(_5512__7_) );
OAI21X1 OAI21X1_1715 ( .gnd(gnd), .vdd(vdd), .A(_1424_), .B(raddr2_0_bF_buf50_), .C(raddr2_1_bF_buf11_), .Y(_4404_) );
AOI21X1 AOI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(regs_20__8_), .B(raddr2_0_bF_buf49_), .C(_4404_), .Y(_4405_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(regs_22__8_), .B(raddr2_0_bF_buf48_), .Y(_4406_) );
OAI21X1 OAI21X1_1716 ( .gnd(gnd), .vdd(vdd), .A(_1326_), .B(raddr2_0_bF_buf47_), .C(_4038__bF_buf2), .Y(_4407_) );
OAI21X1 OAI21X1_1717 ( .gnd(gnd), .vdd(vdd), .A(_4407_), .B(_4406_), .C(_4036__bF_buf3), .Y(_4408_) );
OAI21X1 OAI21X1_1718 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .B(raddr2_0_bF_buf46_), .C(raddr2_1_bF_buf10_), .Y(_4409_) );
AOI21X1 AOI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(regs_16__8_), .B(raddr2_0_bF_buf45_), .C(_4409_), .Y(_4410_) );
NOR2X1 NOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf44_), .B(_1523_), .Y(_4411_) );
NAND2X1 NAND2X1_794 ( .gnd(gnd), .vdd(vdd), .A(regs_18__8_), .B(raddr2_0_bF_buf43_), .Y(_4412_) );
NAND2X1 NAND2X1_795 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf1), .B(_4412_), .Y(_4413_) );
OAI21X1 OAI21X1_1719 ( .gnd(gnd), .vdd(vdd), .A(_4413_), .B(_4411_), .C(raddr2_2_bF_buf10_), .Y(_4414_) );
OAI22X1 OAI22X1_67 ( .gnd(gnd), .vdd(vdd), .A(_4410_), .B(_4414_), .C(_4408_), .D(_4405_), .Y(_4415_) );
NAND2X1 NAND2X1_796 ( .gnd(gnd), .vdd(vdd), .A(regs_28__8_), .B(raddr2_0_bF_buf42_), .Y(_4416_) );
OAI21X1 OAI21X1_1720 ( .gnd(gnd), .vdd(vdd), .A(_2847_), .B(raddr2_0_bF_buf41_), .C(_4416_), .Y(_4417_) );
MUX2X1 MUX2X1_373 ( .gnd(gnd), .vdd(vdd), .A(_4417_), .B(regs_30__8_), .S(raddr2_1_bF_buf9_), .Y(_4418_) );
NAND2X1 NAND2X1_797 ( .gnd(gnd), .vdd(vdd), .A(regs_26__8_), .B(raddr2_0_bF_buf40_), .Y(_4419_) );
OAI21X1 OAI21X1_1721 ( .gnd(gnd), .vdd(vdd), .A(_1159_), .B(raddr2_0_bF_buf39_), .C(_4419_), .Y(_4420_) );
NAND2X1 NAND2X1_798 ( .gnd(gnd), .vdd(vdd), .A(regs_24__8_), .B(raddr2_0_bF_buf38_), .Y(_4421_) );
OAI21X1 OAI21X1_1722 ( .gnd(gnd), .vdd(vdd), .A(_2853_), .B(raddr2_0_bF_buf37_), .C(_4421_), .Y(_4422_) );
MUX2X1 MUX2X1_374 ( .gnd(gnd), .vdd(vdd), .A(_4422_), .B(_4420_), .S(raddr2_1_bF_buf8_), .Y(_4423_) );
MUX2X1 MUX2X1_375 ( .gnd(gnd), .vdd(vdd), .A(_4423_), .B(_4418_), .S(raddr2_2_bF_buf9_), .Y(_4424_) );
MUX2X1 MUX2X1_376 ( .gnd(gnd), .vdd(vdd), .A(_4424_), .B(_4415_), .S(_4033__bF_buf4), .Y(_4425_) );
NAND2X1 NAND2X1_799 ( .gnd(gnd), .vdd(vdd), .A(regs_6__8_), .B(raddr2_0_bF_buf36_), .Y(_4426_) );
OAI21X1 OAI21X1_1723 ( .gnd(gnd), .vdd(vdd), .A(_2117_), .B(raddr2_0_bF_buf35_), .C(_4426_), .Y(_4427_) );
NAND2X1 NAND2X1_800 ( .gnd(gnd), .vdd(vdd), .A(regs_4__8_), .B(raddr2_0_bF_buf34_), .Y(_4428_) );
OAI21X1 OAI21X1_1724 ( .gnd(gnd), .vdd(vdd), .A(_2808_), .B(raddr2_0_bF_buf33_), .C(_4428_), .Y(_4429_) );
MUX2X1 MUX2X1_377 ( .gnd(gnd), .vdd(vdd), .A(_4429_), .B(_4427_), .S(raddr2_1_bF_buf7_), .Y(_4430_) );
NAND2X1 NAND2X1_801 ( .gnd(gnd), .vdd(vdd), .A(regs_2__8_), .B(raddr2_0_bF_buf32_), .Y(_4431_) );
OAI21X1 OAI21X1_1725 ( .gnd(gnd), .vdd(vdd), .A(_2817_), .B(raddr2_0_bF_buf31_), .C(_4431_), .Y(_4432_) );
NAND2X1 NAND2X1_802 ( .gnd(gnd), .vdd(vdd), .A(regs_0__8_), .B(raddr2_0_bF_buf30_), .Y(_4433_) );
OAI21X1 OAI21X1_1726 ( .gnd(gnd), .vdd(vdd), .A(_2814_), .B(raddr2_0_bF_buf29_), .C(_4433_), .Y(_4434_) );
MUX2X1 MUX2X1_378 ( .gnd(gnd), .vdd(vdd), .A(_4434_), .B(_4432_), .S(raddr2_1_bF_buf6_), .Y(_4435_) );
MUX2X1 MUX2X1_379 ( .gnd(gnd), .vdd(vdd), .A(_4435_), .B(_4430_), .S(raddr2_2_bF_buf8_), .Y(_4436_) );
NAND2X1 NAND2X1_803 ( .gnd(gnd), .vdd(vdd), .A(regs_14__8_), .B(raddr2_0_bF_buf28_), .Y(_4437_) );
OAI21X1 OAI21X1_1727 ( .gnd(gnd), .vdd(vdd), .A(_1721_), .B(raddr2_0_bF_buf27_), .C(_4437_), .Y(_4438_) );
NAND2X1 NAND2X1_804 ( .gnd(gnd), .vdd(vdd), .A(regs_12__8_), .B(raddr2_0_bF_buf26_), .Y(_4439_) );
OAI21X1 OAI21X1_1728 ( .gnd(gnd), .vdd(vdd), .A(_1819_), .B(raddr2_0_bF_buf25_), .C(_4439_), .Y(_4440_) );
MUX2X1 MUX2X1_380 ( .gnd(gnd), .vdd(vdd), .A(_4440_), .B(_4438_), .S(raddr2_1_bF_buf5_), .Y(_4441_) );
NAND2X1 NAND2X1_805 ( .gnd(gnd), .vdd(vdd), .A(regs_10__8_), .B(raddr2_0_bF_buf24_), .Y(_4442_) );
OAI21X1 OAI21X1_1729 ( .gnd(gnd), .vdd(vdd), .A(_1918_), .B(raddr2_0_bF_buf23_), .C(_4442_), .Y(_4443_) );
NAND2X1 NAND2X1_806 ( .gnd(gnd), .vdd(vdd), .A(regs_8__8_), .B(raddr2_0_bF_buf22_), .Y(_4444_) );
OAI21X1 OAI21X1_1730 ( .gnd(gnd), .vdd(vdd), .A(_2016_), .B(raddr2_0_bF_buf21_), .C(_4444_), .Y(_4445_) );
MUX2X1 MUX2X1_381 ( .gnd(gnd), .vdd(vdd), .A(_4445_), .B(_4443_), .S(raddr2_1_bF_buf4_), .Y(_4446_) );
MUX2X1 MUX2X1_382 ( .gnd(gnd), .vdd(vdd), .A(_4446_), .B(_4441_), .S(raddr2_2_bF_buf7_), .Y(_4447_) );
MUX2X1 MUX2X1_383 ( .gnd(gnd), .vdd(vdd), .A(_4447_), .B(_4436_), .S(_4033__bF_buf3), .Y(_4448_) );
MUX2X1 MUX2X1_384 ( .gnd(gnd), .vdd(vdd), .A(_4448_), .B(_4425_), .S(raddr2_4_bF_buf1_), .Y(_5512__8_) );
NAND2X1 NAND2X1_807 ( .gnd(gnd), .vdd(vdd), .A(regs_22__9_), .B(raddr2_0_bF_buf20_), .Y(_4449_) );
OAI21X1 OAI21X1_1731 ( .gnd(gnd), .vdd(vdd), .A(_1328_), .B(raddr2_0_bF_buf19_), .C(_4449_), .Y(_4450_) );
NAND2X1 NAND2X1_808 ( .gnd(gnd), .vdd(vdd), .A(regs_20__9_), .B(raddr2_0_bF_buf18_), .Y(_4451_) );
OAI21X1 OAI21X1_1732 ( .gnd(gnd), .vdd(vdd), .A(_1426_), .B(raddr2_0_bF_buf17_), .C(_4451_), .Y(_4452_) );
MUX2X1 MUX2X1_385 ( .gnd(gnd), .vdd(vdd), .A(_4452_), .B(_4450_), .S(raddr2_1_bF_buf3_), .Y(_4453_) );
NAND2X1 NAND2X1_809 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf2), .B(_4453_), .Y(_4454_) );
NAND2X1 NAND2X1_810 ( .gnd(gnd), .vdd(vdd), .A(regs_18__9_), .B(raddr2_0_bF_buf16_), .Y(_4455_) );
OAI21X1 OAI21X1_1733 ( .gnd(gnd), .vdd(vdd), .A(_1525_), .B(raddr2_0_bF_buf15_), .C(_4455_), .Y(_4456_) );
NAND2X1 NAND2X1_811 ( .gnd(gnd), .vdd(vdd), .A(regs_16__9_), .B(raddr2_0_bF_buf14_), .Y(_4457_) );
OAI21X1 OAI21X1_1734 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(raddr2_0_bF_buf13_), .C(_4457_), .Y(_4458_) );
MUX2X1 MUX2X1_386 ( .gnd(gnd), .vdd(vdd), .A(_4458_), .B(_4456_), .S(raddr2_1_bF_buf2_), .Y(_4459_) );
AOI21X1 AOI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(raddr2_2_bF_buf6_), .B(_4459_), .C(_4033__bF_buf2), .Y(_4460_) );
OAI21X1 OAI21X1_1735 ( .gnd(gnd), .vdd(vdd), .A(_1161_), .B(raddr2_0_bF_buf12_), .C(raddr2_2_bF_buf5_), .Y(_4461_) );
AOI21X1 AOI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(regs_26__9_), .B(raddr2_0_bF_buf11_), .C(_4461_), .Y(_4462_) );
OAI21X1 OAI21X1_1736 ( .gnd(gnd), .vdd(vdd), .A(regs_30__9_), .B(raddr2_2_bF_buf4_), .C(_4038__bF_buf0), .Y(_4463_) );
OAI21X1 OAI21X1_1737 ( .gnd(gnd), .vdd(vdd), .A(_2874_), .B(raddr2_0_bF_buf10_), .C(raddr2_2_bF_buf3_), .Y(_4464_) );
AOI21X1 AOI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(regs_24__9_), .B(raddr2_0_bF_buf9_), .C(_4464_), .Y(_4465_) );
NOR2X1 NOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf8_), .B(_2877_), .Y(_4466_) );
NAND2X1 NAND2X1_812 ( .gnd(gnd), .vdd(vdd), .A(regs_28__9_), .B(raddr2_0_bF_buf7_), .Y(_4467_) );
NAND2X1 NAND2X1_813 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf1), .B(_4467_), .Y(_4468_) );
OAI21X1 OAI21X1_1738 ( .gnd(gnd), .vdd(vdd), .A(_4468_), .B(_4466_), .C(raddr2_1_bF_buf1_), .Y(_4469_) );
OAI22X1 OAI22X1_68 ( .gnd(gnd), .vdd(vdd), .A(_4462_), .B(_4463_), .C(_4469_), .D(_4465_), .Y(_4470_) );
AOI22X1 AOI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_4470_), .B(_4033__bF_buf1), .C(_4454_), .D(_4460_), .Y(_4471_) );
OAI21X1 OAI21X1_1739 ( .gnd(gnd), .vdd(vdd), .A(_2886_), .B(raddr2_0_bF_buf6_), .C(raddr2_1_bF_buf0_), .Y(_4472_) );
AOI21X1 AOI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(regs_4__9_), .B(raddr2_0_bF_buf5_), .C(_4472_), .Y(_4473_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(regs_6__9_), .B(raddr2_0_bF_buf4_), .Y(_4474_) );
OAI21X1 OAI21X1_1740 ( .gnd(gnd), .vdd(vdd), .A(_2119_), .B(raddr2_0_bF_buf3_), .C(_4038__bF_buf8), .Y(_4475_) );
OAI21X1 OAI21X1_1741 ( .gnd(gnd), .vdd(vdd), .A(_4475_), .B(_4474_), .C(_4036__bF_buf0), .Y(_4476_) );
OAI21X1 OAI21X1_1742 ( .gnd(gnd), .vdd(vdd), .A(_2893_), .B(raddr2_0_bF_buf2_), .C(raddr2_1_bF_buf14_bF_buf2_), .Y(_4477_) );
AOI21X1 AOI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(regs_0__9_), .B(raddr2_0_bF_buf1_), .C(_4477_), .Y(_4478_) );
NOR2X1 NOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf0_), .B(_2890_), .Y(_4479_) );
NAND2X1 NAND2X1_814 ( .gnd(gnd), .vdd(vdd), .A(regs_2__9_), .B(raddr2_0_bF_buf96_), .Y(_4480_) );
NAND2X1 NAND2X1_815 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf7), .B(_4480_), .Y(_4481_) );
OAI21X1 OAI21X1_1743 ( .gnd(gnd), .vdd(vdd), .A(_4481_), .B(_4479_), .C(raddr2_2_bF_buf2_), .Y(_4482_) );
OAI22X1 OAI22X1_69 ( .gnd(gnd), .vdd(vdd), .A(_4478_), .B(_4482_), .C(_4476_), .D(_4473_), .Y(_4483_) );
NAND2X1 NAND2X1_816 ( .gnd(gnd), .vdd(vdd), .A(regs_10__9_), .B(raddr2_0_bF_buf95_), .Y(_4484_) );
OAI21X1 OAI21X1_1744 ( .gnd(gnd), .vdd(vdd), .A(_1920_), .B(raddr2_0_bF_buf94_), .C(_4484_), .Y(_4485_) );
NAND2X1 NAND2X1_817 ( .gnd(gnd), .vdd(vdd), .A(regs_8__9_), .B(raddr2_0_bF_buf93_), .Y(_4486_) );
OAI21X1 OAI21X1_1745 ( .gnd(gnd), .vdd(vdd), .A(_2018_), .B(raddr2_0_bF_buf92_), .C(_4486_), .Y(_4487_) );
MUX2X1 MUX2X1_387 ( .gnd(gnd), .vdd(vdd), .A(_4487_), .B(_4485_), .S(raddr2_1_bF_buf13_bF_buf2_), .Y(_4488_) );
NAND2X1 NAND2X1_818 ( .gnd(gnd), .vdd(vdd), .A(regs_14__9_), .B(raddr2_0_bF_buf91_), .Y(_4489_) );
OAI21X1 OAI21X1_1746 ( .gnd(gnd), .vdd(vdd), .A(_1723_), .B(raddr2_0_bF_buf90_), .C(_4489_), .Y(_4490_) );
NAND2X1 NAND2X1_819 ( .gnd(gnd), .vdd(vdd), .A(regs_12__9_), .B(raddr2_0_bF_buf89_), .Y(_4491_) );
OAI21X1 OAI21X1_1747 ( .gnd(gnd), .vdd(vdd), .A(_1821_), .B(raddr2_0_bF_buf88_), .C(_4491_), .Y(_4492_) );
MUX2X1 MUX2X1_388 ( .gnd(gnd), .vdd(vdd), .A(_4492_), .B(_4490_), .S(raddr2_1_bF_buf12_bF_buf2_), .Y(_4493_) );
MUX2X1 MUX2X1_389 ( .gnd(gnd), .vdd(vdd), .A(_4493_), .B(_4488_), .S(_4036__bF_buf8), .Y(_4494_) );
MUX2X1 MUX2X1_390 ( .gnd(gnd), .vdd(vdd), .A(_4494_), .B(_4483_), .S(_4033__bF_buf0), .Y(_4495_) );
MUX2X1 MUX2X1_391 ( .gnd(gnd), .vdd(vdd), .A(_4495_), .B(_4471_), .S(raddr2_4_bF_buf0_), .Y(_5512__9_) );
OAI21X1 OAI21X1_1748 ( .gnd(gnd), .vdd(vdd), .A(_2935_), .B(raddr2_0_bF_buf87_), .C(raddr2_1_bF_buf11_), .Y(_4496_) );
AOI21X1 AOI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(regs_4__10_), .B(raddr2_0_bF_buf86_), .C(_4496_), .Y(_4497_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(regs_6__10_), .B(raddr2_0_bF_buf85_), .Y(_4498_) );
OAI21X1 OAI21X1_1749 ( .gnd(gnd), .vdd(vdd), .A(_2121_), .B(raddr2_0_bF_buf84_), .C(_4038__bF_buf6), .Y(_4499_) );
OAI21X1 OAI21X1_1750 ( .gnd(gnd), .vdd(vdd), .A(_4499_), .B(_4498_), .C(_4036__bF_buf7), .Y(_4500_) );
OAI21X1 OAI21X1_1751 ( .gnd(gnd), .vdd(vdd), .A(_2941_), .B(raddr2_0_bF_buf83_), .C(raddr2_1_bF_buf10_), .Y(_4501_) );
AOI21X1 AOI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(regs_0__10_), .B(raddr2_0_bF_buf82_), .C(_4501_), .Y(_4502_) );
NOR2X1 NOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf81_), .B(_2944_), .Y(_4503_) );
NAND2X1 NAND2X1_820 ( .gnd(gnd), .vdd(vdd), .A(regs_2__10_), .B(raddr2_0_bF_buf80_), .Y(_4504_) );
NAND2X1 NAND2X1_821 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf5), .B(_4504_), .Y(_4505_) );
OAI21X1 OAI21X1_1752 ( .gnd(gnd), .vdd(vdd), .A(_4505_), .B(_4503_), .C(raddr2_2_bF_buf1_), .Y(_4506_) );
OAI22X1 OAI22X1_70 ( .gnd(gnd), .vdd(vdd), .A(_4502_), .B(_4506_), .C(_4500_), .D(_4497_), .Y(_4507_) );
NAND2X1 NAND2X1_822 ( .gnd(gnd), .vdd(vdd), .A(regs_10__10_), .B(raddr2_0_bF_buf79_), .Y(_4508_) );
OAI21X1 OAI21X1_1753 ( .gnd(gnd), .vdd(vdd), .A(_1922_), .B(raddr2_0_bF_buf78_), .C(_4508_), .Y(_4509_) );
NAND2X1 NAND2X1_823 ( .gnd(gnd), .vdd(vdd), .A(regs_8__10_), .B(raddr2_0_bF_buf77_), .Y(_4510_) );
OAI21X1 OAI21X1_1754 ( .gnd(gnd), .vdd(vdd), .A(_2020_), .B(raddr2_0_bF_buf76_), .C(_4510_), .Y(_4511_) );
MUX2X1 MUX2X1_392 ( .gnd(gnd), .vdd(vdd), .A(_4511_), .B(_4509_), .S(raddr2_1_bF_buf9_), .Y(_4512_) );
NAND2X1 NAND2X1_824 ( .gnd(gnd), .vdd(vdd), .A(regs_14__10_), .B(raddr2_0_bF_buf75_), .Y(_4513_) );
OAI21X1 OAI21X1_1755 ( .gnd(gnd), .vdd(vdd), .A(_1725_), .B(raddr2_0_bF_buf74_), .C(_4513_), .Y(_4514_) );
NAND2X1 NAND2X1_825 ( .gnd(gnd), .vdd(vdd), .A(regs_12__10_), .B(raddr2_0_bF_buf73_), .Y(_4515_) );
OAI21X1 OAI21X1_1756 ( .gnd(gnd), .vdd(vdd), .A(_1823_), .B(raddr2_0_bF_buf72_), .C(_4515_), .Y(_4516_) );
MUX2X1 MUX2X1_393 ( .gnd(gnd), .vdd(vdd), .A(_4516_), .B(_4514_), .S(raddr2_1_bF_buf8_), .Y(_4517_) );
MUX2X1 MUX2X1_394 ( .gnd(gnd), .vdd(vdd), .A(_4517_), .B(_4512_), .S(_4036__bF_buf6), .Y(_4518_) );
MUX2X1 MUX2X1_395 ( .gnd(gnd), .vdd(vdd), .A(_4518_), .B(_4507_), .S(_4033__bF_buf7), .Y(_4519_) );
OAI21X1 OAI21X1_1757 ( .gnd(gnd), .vdd(vdd), .A(_1625_), .B(raddr2_0_bF_buf71_), .C(raddr2_1_bF_buf7_), .Y(_4520_) );
AOI21X1 AOI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(regs_16__10_), .B(raddr2_0_bF_buf70_), .C(_4520_), .Y(_4521_) );
NOR2X1 NOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf69_), .B(_1527_), .Y(_4522_) );
NAND2X1 NAND2X1_826 ( .gnd(gnd), .vdd(vdd), .A(regs_18__10_), .B(raddr2_0_bF_buf68_), .Y(_4523_) );
NAND2X1 NAND2X1_827 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf4), .B(_4523_), .Y(_4524_) );
OAI21X1 OAI21X1_1758 ( .gnd(gnd), .vdd(vdd), .A(_4524_), .B(_4522_), .C(raddr2_2_bF_buf0_), .Y(_4525_) );
OAI21X1 OAI21X1_1759 ( .gnd(gnd), .vdd(vdd), .A(_1428_), .B(raddr2_0_bF_buf67_), .C(raddr2_1_bF_buf6_), .Y(_4526_) );
AOI21X1 AOI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(regs_20__10_), .B(raddr2_0_bF_buf66_), .C(_4526_), .Y(_4527_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(regs_22__10_), .B(raddr2_0_bF_buf65_), .Y(_4528_) );
OAI21X1 OAI21X1_1760 ( .gnd(gnd), .vdd(vdd), .A(_1330_), .B(raddr2_0_bF_buf64_), .C(_4038__bF_buf3), .Y(_4529_) );
OAI21X1 OAI21X1_1761 ( .gnd(gnd), .vdd(vdd), .A(_4529_), .B(_4528_), .C(_4036__bF_buf5), .Y(_4530_) );
OAI22X1 OAI22X1_71 ( .gnd(gnd), .vdd(vdd), .A(_4521_), .B(_4525_), .C(_4530_), .D(_4527_), .Y(_4531_) );
NAND2X1 NAND2X1_828 ( .gnd(gnd), .vdd(vdd), .A(regs_28__10_), .B(raddr2_0_bF_buf63_), .Y(_4532_) );
OAI21X1 OAI21X1_1762 ( .gnd(gnd), .vdd(vdd), .A(_2928_), .B(raddr2_0_bF_buf62_), .C(_4532_), .Y(_4533_) );
MUX2X1 MUX2X1_396 ( .gnd(gnd), .vdd(vdd), .A(_4533_), .B(regs_30__10_), .S(raddr2_1_bF_buf5_), .Y(_4534_) );
NAND2X1 NAND2X1_829 ( .gnd(gnd), .vdd(vdd), .A(regs_26__10_), .B(raddr2_0_bF_buf61_), .Y(_4535_) );
OAI21X1 OAI21X1_1763 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(raddr2_0_bF_buf60_), .C(_4535_), .Y(_4536_) );
NAND2X1 NAND2X1_830 ( .gnd(gnd), .vdd(vdd), .A(regs_24__10_), .B(raddr2_0_bF_buf59_), .Y(_4537_) );
OAI21X1 OAI21X1_1764 ( .gnd(gnd), .vdd(vdd), .A(_2925_), .B(raddr2_0_bF_buf58_), .C(_4537_), .Y(_4538_) );
MUX2X1 MUX2X1_397 ( .gnd(gnd), .vdd(vdd), .A(_4538_), .B(_4536_), .S(raddr2_1_bF_buf4_), .Y(_4539_) );
MUX2X1 MUX2X1_398 ( .gnd(gnd), .vdd(vdd), .A(_4539_), .B(_4534_), .S(raddr2_2_bF_buf10_), .Y(_4540_) );
MUX2X1 MUX2X1_399 ( .gnd(gnd), .vdd(vdd), .A(_4540_), .B(_4531_), .S(_4033__bF_buf6), .Y(_4541_) );
MUX2X1 MUX2X1_400 ( .gnd(gnd), .vdd(vdd), .A(_4519_), .B(_4541_), .S(raddr2_4_bF_buf4_), .Y(_5512__10_) );
OAI21X1 OAI21X1_1765 ( .gnd(gnd), .vdd(vdd), .A(_2962_), .B(raddr2_0_bF_buf57_), .C(raddr2_1_bF_buf3_), .Y(_4542_) );
AOI21X1 AOI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(regs_4__11_), .B(raddr2_0_bF_buf56_), .C(_4542_), .Y(_4543_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(regs_6__11_), .B(raddr2_0_bF_buf55_), .Y(_4544_) );
OAI21X1 OAI21X1_1766 ( .gnd(gnd), .vdd(vdd), .A(_2123_), .B(raddr2_0_bF_buf54_), .C(_4038__bF_buf2), .Y(_4545_) );
OAI21X1 OAI21X1_1767 ( .gnd(gnd), .vdd(vdd), .A(_4545_), .B(_4544_), .C(_4036__bF_buf4), .Y(_4546_) );
OAI21X1 OAI21X1_1768 ( .gnd(gnd), .vdd(vdd), .A(_2968_), .B(raddr2_0_bF_buf53_), .C(raddr2_1_bF_buf2_), .Y(_4547_) );
AOI21X1 AOI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(regs_0__11_), .B(raddr2_0_bF_buf52_), .C(_4547_), .Y(_4548_) );
NOR2X1 NOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf51_), .B(_2971_), .Y(_4549_) );
NAND2X1 NAND2X1_831 ( .gnd(gnd), .vdd(vdd), .A(regs_2__11_), .B(raddr2_0_bF_buf50_), .Y(_4550_) );
NAND2X1 NAND2X1_832 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf1), .B(_4550_), .Y(_4551_) );
OAI21X1 OAI21X1_1769 ( .gnd(gnd), .vdd(vdd), .A(_4551_), .B(_4549_), .C(raddr2_2_bF_buf9_), .Y(_4552_) );
OAI22X1 OAI22X1_72 ( .gnd(gnd), .vdd(vdd), .A(_4548_), .B(_4552_), .C(_4546_), .D(_4543_), .Y(_4553_) );
NAND2X1 NAND2X1_833 ( .gnd(gnd), .vdd(vdd), .A(regs_10__11_), .B(raddr2_0_bF_buf49_), .Y(_4554_) );
OAI21X1 OAI21X1_1770 ( .gnd(gnd), .vdd(vdd), .A(_1924_), .B(raddr2_0_bF_buf48_), .C(_4554_), .Y(_4555_) );
NAND2X1 NAND2X1_834 ( .gnd(gnd), .vdd(vdd), .A(regs_8__11_), .B(raddr2_0_bF_buf47_), .Y(_4556_) );
OAI21X1 OAI21X1_1771 ( .gnd(gnd), .vdd(vdd), .A(_2022_), .B(raddr2_0_bF_buf46_), .C(_4556_), .Y(_4557_) );
MUX2X1 MUX2X1_401 ( .gnd(gnd), .vdd(vdd), .A(_4557_), .B(_4555_), .S(raddr2_1_bF_buf1_), .Y(_4558_) );
NAND2X1 NAND2X1_835 ( .gnd(gnd), .vdd(vdd), .A(regs_14__11_), .B(raddr2_0_bF_buf45_), .Y(_4559_) );
OAI21X1 OAI21X1_1772 ( .gnd(gnd), .vdd(vdd), .A(_1727_), .B(raddr2_0_bF_buf44_), .C(_4559_), .Y(_4560_) );
NAND2X1 NAND2X1_836 ( .gnd(gnd), .vdd(vdd), .A(regs_12__11_), .B(raddr2_0_bF_buf43_), .Y(_4561_) );
OAI21X1 OAI21X1_1773 ( .gnd(gnd), .vdd(vdd), .A(_1825_), .B(raddr2_0_bF_buf42_), .C(_4561_), .Y(_4562_) );
MUX2X1 MUX2X1_402 ( .gnd(gnd), .vdd(vdd), .A(_4562_), .B(_4560_), .S(raddr2_1_bF_buf0_), .Y(_4563_) );
MUX2X1 MUX2X1_403 ( .gnd(gnd), .vdd(vdd), .A(_4563_), .B(_4558_), .S(_4036__bF_buf3), .Y(_4564_) );
MUX2X1 MUX2X1_404 ( .gnd(gnd), .vdd(vdd), .A(_4564_), .B(_4553_), .S(_4033__bF_buf5), .Y(_4565_) );
OAI21X1 OAI21X1_1774 ( .gnd(gnd), .vdd(vdd), .A(_1627_), .B(raddr2_0_bF_buf41_), .C(raddr2_1_bF_buf14_bF_buf1_), .Y(_4566_) );
AOI21X1 AOI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(regs_16__11_), .B(raddr2_0_bF_buf40_), .C(_4566_), .Y(_4567_) );
NOR2X1 NOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf39_), .B(_1529_), .Y(_4568_) );
NAND2X1 NAND2X1_837 ( .gnd(gnd), .vdd(vdd), .A(regs_18__11_), .B(raddr2_0_bF_buf38_), .Y(_4569_) );
NAND2X1 NAND2X1_838 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf0), .B(_4569_), .Y(_4570_) );
OAI21X1 OAI21X1_1775 ( .gnd(gnd), .vdd(vdd), .A(_4570_), .B(_4568_), .C(raddr2_2_bF_buf8_), .Y(_4571_) );
OAI21X1 OAI21X1_1776 ( .gnd(gnd), .vdd(vdd), .A(_1430_), .B(raddr2_0_bF_buf37_), .C(raddr2_1_bF_buf13_bF_buf1_), .Y(_4572_) );
AOI21X1 AOI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(regs_20__11_), .B(raddr2_0_bF_buf36_), .C(_4572_), .Y(_4573_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(regs_22__11_), .B(raddr2_0_bF_buf35_), .Y(_4574_) );
OAI21X1 OAI21X1_1777 ( .gnd(gnd), .vdd(vdd), .A(_1332_), .B(raddr2_0_bF_buf34_), .C(_4038__bF_buf8), .Y(_4575_) );
OAI21X1 OAI21X1_1778 ( .gnd(gnd), .vdd(vdd), .A(_4575_), .B(_4574_), .C(_4036__bF_buf2), .Y(_4576_) );
OAI22X1 OAI22X1_73 ( .gnd(gnd), .vdd(vdd), .A(_4567_), .B(_4571_), .C(_4576_), .D(_4573_), .Y(_4577_) );
NAND2X1 NAND2X1_839 ( .gnd(gnd), .vdd(vdd), .A(regs_28__11_), .B(raddr2_0_bF_buf33_), .Y(_4578_) );
OAI21X1 OAI21X1_1779 ( .gnd(gnd), .vdd(vdd), .A(_3001_), .B(raddr2_0_bF_buf32_), .C(_4578_), .Y(_4579_) );
MUX2X1 MUX2X1_405 ( .gnd(gnd), .vdd(vdd), .A(_4579_), .B(regs_30__11_), .S(raddr2_1_bF_buf12_bF_buf1_), .Y(_4580_) );
NAND2X1 NAND2X1_840 ( .gnd(gnd), .vdd(vdd), .A(regs_26__11_), .B(raddr2_0_bF_buf31_), .Y(_4581_) );
OAI21X1 OAI21X1_1780 ( .gnd(gnd), .vdd(vdd), .A(_1165_), .B(raddr2_0_bF_buf30_), .C(_4581_), .Y(_4582_) );
NAND2X1 NAND2X1_841 ( .gnd(gnd), .vdd(vdd), .A(regs_24__11_), .B(raddr2_0_bF_buf29_), .Y(_4583_) );
OAI21X1 OAI21X1_1781 ( .gnd(gnd), .vdd(vdd), .A(_3007_), .B(raddr2_0_bF_buf28_), .C(_4583_), .Y(_4584_) );
MUX2X1 MUX2X1_406 ( .gnd(gnd), .vdd(vdd), .A(_4584_), .B(_4582_), .S(raddr2_1_bF_buf11_), .Y(_4585_) );
MUX2X1 MUX2X1_407 ( .gnd(gnd), .vdd(vdd), .A(_4585_), .B(_4580_), .S(raddr2_2_bF_buf7_), .Y(_4586_) );
MUX2X1 MUX2X1_408 ( .gnd(gnd), .vdd(vdd), .A(_4586_), .B(_4577_), .S(_4033__bF_buf4), .Y(_4587_) );
MUX2X1 MUX2X1_409 ( .gnd(gnd), .vdd(vdd), .A(_4565_), .B(_4587_), .S(raddr2_4_bF_buf3_), .Y(_5512__11_) );
OAI21X1 OAI21X1_1782 ( .gnd(gnd), .vdd(vdd), .A(_3013_), .B(raddr2_0_bF_buf27_), .C(raddr2_1_bF_buf10_), .Y(_4588_) );
AOI21X1 AOI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(regs_4__12_), .B(raddr2_0_bF_buf26_), .C(_4588_), .Y(_4589_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(regs_6__12_), .B(raddr2_0_bF_buf25_), .Y(_4590_) );
OAI21X1 OAI21X1_1783 ( .gnd(gnd), .vdd(vdd), .A(_2125_), .B(raddr2_0_bF_buf24_), .C(_4038__bF_buf7), .Y(_4591_) );
OAI21X1 OAI21X1_1784 ( .gnd(gnd), .vdd(vdd), .A(_4591_), .B(_4590_), .C(_4036__bF_buf1), .Y(_4592_) );
OAI21X1 OAI21X1_1785 ( .gnd(gnd), .vdd(vdd), .A(_3019_), .B(raddr2_0_bF_buf23_), .C(raddr2_1_bF_buf9_), .Y(_4593_) );
AOI21X1 AOI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(regs_0__12_), .B(raddr2_0_bF_buf22_), .C(_4593_), .Y(_4594_) );
NOR2X1 NOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf21_), .B(_3022_), .Y(_4595_) );
NAND2X1 NAND2X1_842 ( .gnd(gnd), .vdd(vdd), .A(regs_2__12_), .B(raddr2_0_bF_buf20_), .Y(_4596_) );
NAND2X1 NAND2X1_843 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf6), .B(_4596_), .Y(_4597_) );
OAI21X1 OAI21X1_1786 ( .gnd(gnd), .vdd(vdd), .A(_4597_), .B(_4595_), .C(raddr2_2_bF_buf6_), .Y(_4598_) );
OAI22X1 OAI22X1_74 ( .gnd(gnd), .vdd(vdd), .A(_4594_), .B(_4598_), .C(_4592_), .D(_4589_), .Y(_4599_) );
NAND2X1 NAND2X1_844 ( .gnd(gnd), .vdd(vdd), .A(regs_10__12_), .B(raddr2_0_bF_buf19_), .Y(_4600_) );
OAI21X1 OAI21X1_1787 ( .gnd(gnd), .vdd(vdd), .A(_1926_), .B(raddr2_0_bF_buf18_), .C(_4600_), .Y(_4601_) );
NAND2X1 NAND2X1_845 ( .gnd(gnd), .vdd(vdd), .A(regs_8__12_), .B(raddr2_0_bF_buf17_), .Y(_4602_) );
OAI21X1 OAI21X1_1788 ( .gnd(gnd), .vdd(vdd), .A(_2024_), .B(raddr2_0_bF_buf16_), .C(_4602_), .Y(_4603_) );
MUX2X1 MUX2X1_410 ( .gnd(gnd), .vdd(vdd), .A(_4603_), .B(_4601_), .S(raddr2_1_bF_buf8_), .Y(_4604_) );
NAND2X1 NAND2X1_846 ( .gnd(gnd), .vdd(vdd), .A(regs_14__12_), .B(raddr2_0_bF_buf15_), .Y(_4605_) );
OAI21X1 OAI21X1_1789 ( .gnd(gnd), .vdd(vdd), .A(_1729_), .B(raddr2_0_bF_buf14_), .C(_4605_), .Y(_4606_) );
NAND2X1 NAND2X1_847 ( .gnd(gnd), .vdd(vdd), .A(regs_12__12_), .B(raddr2_0_bF_buf13_), .Y(_4607_) );
OAI21X1 OAI21X1_1790 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .B(raddr2_0_bF_buf12_), .C(_4607_), .Y(_4608_) );
MUX2X1 MUX2X1_411 ( .gnd(gnd), .vdd(vdd), .A(_4608_), .B(_4606_), .S(raddr2_1_bF_buf7_), .Y(_4609_) );
MUX2X1 MUX2X1_412 ( .gnd(gnd), .vdd(vdd), .A(_4609_), .B(_4604_), .S(_4036__bF_buf0), .Y(_4610_) );
MUX2X1 MUX2X1_413 ( .gnd(gnd), .vdd(vdd), .A(_4610_), .B(_4599_), .S(_4033__bF_buf3), .Y(_4611_) );
OAI21X1 OAI21X1_1791 ( .gnd(gnd), .vdd(vdd), .A(_1629_), .B(raddr2_0_bF_buf11_), .C(raddr2_1_bF_buf6_), .Y(_4612_) );
AOI21X1 AOI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(regs_16__12_), .B(raddr2_0_bF_buf10_), .C(_4612_), .Y(_4613_) );
NOR2X1 NOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf9_), .B(_1531_), .Y(_4614_) );
NAND2X1 NAND2X1_848 ( .gnd(gnd), .vdd(vdd), .A(regs_18__12_), .B(raddr2_0_bF_buf8_), .Y(_4615_) );
NAND2X1 NAND2X1_849 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf5), .B(_4615_), .Y(_4616_) );
OAI21X1 OAI21X1_1792 ( .gnd(gnd), .vdd(vdd), .A(_4616_), .B(_4614_), .C(raddr2_2_bF_buf5_), .Y(_4617_) );
OAI21X1 OAI21X1_1793 ( .gnd(gnd), .vdd(vdd), .A(_1432_), .B(raddr2_0_bF_buf7_), .C(raddr2_1_bF_buf5_), .Y(_4618_) );
AOI21X1 AOI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(regs_20__12_), .B(raddr2_0_bF_buf6_), .C(_4618_), .Y(_4619_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(regs_22__12_), .B(raddr2_0_bF_buf5_), .Y(_4620_) );
OAI21X1 OAI21X1_1794 ( .gnd(gnd), .vdd(vdd), .A(_1334_), .B(raddr2_0_bF_buf4_), .C(_4038__bF_buf4), .Y(_4621_) );
OAI21X1 OAI21X1_1795 ( .gnd(gnd), .vdd(vdd), .A(_4621_), .B(_4620_), .C(_4036__bF_buf8), .Y(_4622_) );
OAI22X1 OAI22X1_75 ( .gnd(gnd), .vdd(vdd), .A(_4613_), .B(_4617_), .C(_4622_), .D(_4619_), .Y(_4623_) );
NAND2X1 NAND2X1_850 ( .gnd(gnd), .vdd(vdd), .A(regs_28__12_), .B(raddr2_0_bF_buf3_), .Y(_4624_) );
OAI21X1 OAI21X1_1796 ( .gnd(gnd), .vdd(vdd), .A(_3052_), .B(raddr2_0_bF_buf2_), .C(_4624_), .Y(_4625_) );
MUX2X1 MUX2X1_414 ( .gnd(gnd), .vdd(vdd), .A(_4625_), .B(regs_30__12_), .S(raddr2_1_bF_buf4_), .Y(_4626_) );
NAND2X1 NAND2X1_851 ( .gnd(gnd), .vdd(vdd), .A(regs_26__12_), .B(raddr2_0_bF_buf1_), .Y(_4627_) );
OAI21X1 OAI21X1_1797 ( .gnd(gnd), .vdd(vdd), .A(_1167_), .B(raddr2_0_bF_buf0_), .C(_4627_), .Y(_4628_) );
NAND2X1 NAND2X1_852 ( .gnd(gnd), .vdd(vdd), .A(regs_24__12_), .B(raddr2_0_bF_buf96_), .Y(_4629_) );
OAI21X1 OAI21X1_1798 ( .gnd(gnd), .vdd(vdd), .A(_3058_), .B(raddr2_0_bF_buf95_), .C(_4629_), .Y(_4630_) );
MUX2X1 MUX2X1_415 ( .gnd(gnd), .vdd(vdd), .A(_4630_), .B(_4628_), .S(raddr2_1_bF_buf3_), .Y(_4631_) );
MUX2X1 MUX2X1_416 ( .gnd(gnd), .vdd(vdd), .A(_4631_), .B(_4626_), .S(raddr2_2_bF_buf4_), .Y(_4632_) );
MUX2X1 MUX2X1_417 ( .gnd(gnd), .vdd(vdd), .A(_4632_), .B(_4623_), .S(_4033__bF_buf2), .Y(_4633_) );
MUX2X1 MUX2X1_418 ( .gnd(gnd), .vdd(vdd), .A(_4611_), .B(_4633_), .S(raddr2_4_bF_buf2_), .Y(_5512__12_) );
OAI21X1 OAI21X1_1799 ( .gnd(gnd), .vdd(vdd), .A(_3064_), .B(raddr2_0_bF_buf94_), .C(raddr2_1_bF_buf2_), .Y(_4634_) );
AOI21X1 AOI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(regs_4__13_), .B(raddr2_0_bF_buf93_), .C(_4634_), .Y(_4635_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(regs_6__13_), .B(raddr2_0_bF_buf92_), .Y(_4636_) );
OAI21X1 OAI21X1_1800 ( .gnd(gnd), .vdd(vdd), .A(_2127_), .B(raddr2_0_bF_buf91_), .C(_4038__bF_buf3), .Y(_4637_) );
OAI21X1 OAI21X1_1801 ( .gnd(gnd), .vdd(vdd), .A(_4637_), .B(_4636_), .C(_4036__bF_buf7), .Y(_4638_) );
OAI21X1 OAI21X1_1802 ( .gnd(gnd), .vdd(vdd), .A(_3070_), .B(raddr2_0_bF_buf90_), .C(raddr2_1_bF_buf1_), .Y(_4639_) );
AOI21X1 AOI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(regs_0__13_), .B(raddr2_0_bF_buf89_), .C(_4639_), .Y(_4640_) );
NOR2X1 NOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf88_), .B(_3073_), .Y(_4641_) );
NAND2X1 NAND2X1_853 ( .gnd(gnd), .vdd(vdd), .A(regs_2__13_), .B(raddr2_0_bF_buf87_), .Y(_4642_) );
NAND2X1 NAND2X1_854 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf2), .B(_4642_), .Y(_4643_) );
OAI21X1 OAI21X1_1803 ( .gnd(gnd), .vdd(vdd), .A(_4643_), .B(_4641_), .C(raddr2_2_bF_buf3_), .Y(_4644_) );
OAI22X1 OAI22X1_76 ( .gnd(gnd), .vdd(vdd), .A(_4640_), .B(_4644_), .C(_4638_), .D(_4635_), .Y(_4645_) );
NAND2X1 NAND2X1_855 ( .gnd(gnd), .vdd(vdd), .A(regs_10__13_), .B(raddr2_0_bF_buf86_), .Y(_4646_) );
OAI21X1 OAI21X1_1804 ( .gnd(gnd), .vdd(vdd), .A(_1928_), .B(raddr2_0_bF_buf85_), .C(_4646_), .Y(_4647_) );
NAND2X1 NAND2X1_856 ( .gnd(gnd), .vdd(vdd), .A(regs_8__13_), .B(raddr2_0_bF_buf84_), .Y(_4648_) );
OAI21X1 OAI21X1_1805 ( .gnd(gnd), .vdd(vdd), .A(_2026_), .B(raddr2_0_bF_buf83_), .C(_4648_), .Y(_4649_) );
MUX2X1 MUX2X1_419 ( .gnd(gnd), .vdd(vdd), .A(_4649_), .B(_4647_), .S(raddr2_1_bF_buf0_), .Y(_4650_) );
NAND2X1 NAND2X1_857 ( .gnd(gnd), .vdd(vdd), .A(regs_14__13_), .B(raddr2_0_bF_buf82_), .Y(_4651_) );
OAI21X1 OAI21X1_1806 ( .gnd(gnd), .vdd(vdd), .A(_1731_), .B(raddr2_0_bF_buf81_), .C(_4651_), .Y(_4652_) );
NAND2X1 NAND2X1_858 ( .gnd(gnd), .vdd(vdd), .A(regs_12__13_), .B(raddr2_0_bF_buf80_), .Y(_4653_) );
OAI21X1 OAI21X1_1807 ( .gnd(gnd), .vdd(vdd), .A(_1829_), .B(raddr2_0_bF_buf79_), .C(_4653_), .Y(_4654_) );
MUX2X1 MUX2X1_420 ( .gnd(gnd), .vdd(vdd), .A(_4654_), .B(_4652_), .S(raddr2_1_bF_buf14_bF_buf0_), .Y(_4655_) );
MUX2X1 MUX2X1_421 ( .gnd(gnd), .vdd(vdd), .A(_4655_), .B(_4650_), .S(_4036__bF_buf6), .Y(_4656_) );
MUX2X1 MUX2X1_422 ( .gnd(gnd), .vdd(vdd), .A(_4656_), .B(_4645_), .S(_4033__bF_buf1), .Y(_4657_) );
OAI21X1 OAI21X1_1808 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .B(raddr2_0_bF_buf78_), .C(raddr2_1_bF_buf13_bF_buf0_), .Y(_4658_) );
AOI21X1 AOI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(regs_16__13_), .B(raddr2_0_bF_buf77_), .C(_4658_), .Y(_4659_) );
NOR2X1 NOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf76_), .B(_1533_), .Y(_4660_) );
NAND2X1 NAND2X1_859 ( .gnd(gnd), .vdd(vdd), .A(regs_18__13_), .B(raddr2_0_bF_buf75_), .Y(_4661_) );
NAND2X1 NAND2X1_860 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf1), .B(_4661_), .Y(_4662_) );
OAI21X1 OAI21X1_1809 ( .gnd(gnd), .vdd(vdd), .A(_4662_), .B(_4660_), .C(raddr2_2_bF_buf2_), .Y(_4663_) );
OAI21X1 OAI21X1_1810 ( .gnd(gnd), .vdd(vdd), .A(_1434_), .B(raddr2_0_bF_buf74_), .C(raddr2_1_bF_buf12_bF_buf0_), .Y(_4664_) );
AOI21X1 AOI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(regs_20__13_), .B(raddr2_0_bF_buf73_), .C(_4664_), .Y(_4665_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(regs_22__13_), .B(raddr2_0_bF_buf72_), .Y(_4666_) );
OAI21X1 OAI21X1_1811 ( .gnd(gnd), .vdd(vdd), .A(_1336_), .B(raddr2_0_bF_buf71_), .C(_4038__bF_buf0), .Y(_4667_) );
OAI21X1 OAI21X1_1812 ( .gnd(gnd), .vdd(vdd), .A(_4667_), .B(_4666_), .C(_4036__bF_buf5), .Y(_4668_) );
OAI22X1 OAI22X1_77 ( .gnd(gnd), .vdd(vdd), .A(_4659_), .B(_4663_), .C(_4668_), .D(_4665_), .Y(_4669_) );
NAND2X1 NAND2X1_861 ( .gnd(gnd), .vdd(vdd), .A(regs_28__13_), .B(raddr2_0_bF_buf70_), .Y(_4670_) );
OAI21X1 OAI21X1_1813 ( .gnd(gnd), .vdd(vdd), .A(_3103_), .B(raddr2_0_bF_buf69_), .C(_4670_), .Y(_4671_) );
MUX2X1 MUX2X1_423 ( .gnd(gnd), .vdd(vdd), .A(_4671_), .B(regs_30__13_), .S(raddr2_1_bF_buf11_), .Y(_4672_) );
NAND2X1 NAND2X1_862 ( .gnd(gnd), .vdd(vdd), .A(regs_26__13_), .B(raddr2_0_bF_buf68_), .Y(_4673_) );
OAI21X1 OAI21X1_1814 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(raddr2_0_bF_buf67_), .C(_4673_), .Y(_4674_) );
NAND2X1 NAND2X1_863 ( .gnd(gnd), .vdd(vdd), .A(regs_24__13_), .B(raddr2_0_bF_buf66_), .Y(_4675_) );
OAI21X1 OAI21X1_1815 ( .gnd(gnd), .vdd(vdd), .A(_3109_), .B(raddr2_0_bF_buf65_), .C(_4675_), .Y(_4676_) );
MUX2X1 MUX2X1_424 ( .gnd(gnd), .vdd(vdd), .A(_4676_), .B(_4674_), .S(raddr2_1_bF_buf10_), .Y(_4677_) );
MUX2X1 MUX2X1_425 ( .gnd(gnd), .vdd(vdd), .A(_4677_), .B(_4672_), .S(raddr2_2_bF_buf1_), .Y(_4678_) );
MUX2X1 MUX2X1_426 ( .gnd(gnd), .vdd(vdd), .A(_4678_), .B(_4669_), .S(_4033__bF_buf0), .Y(_4679_) );
MUX2X1 MUX2X1_427 ( .gnd(gnd), .vdd(vdd), .A(_4657_), .B(_4679_), .S(raddr2_4_bF_buf1_), .Y(_5512__13_) );
NAND2X1 NAND2X1_864 ( .gnd(gnd), .vdd(vdd), .A(regs_22__14_), .B(raddr2_0_bF_buf64_), .Y(_4680_) );
OAI21X1 OAI21X1_1816 ( .gnd(gnd), .vdd(vdd), .A(_1338_), .B(raddr2_0_bF_buf63_), .C(_4680_), .Y(_4681_) );
NAND2X1 NAND2X1_865 ( .gnd(gnd), .vdd(vdd), .A(regs_20__14_), .B(raddr2_0_bF_buf62_), .Y(_4682_) );
OAI21X1 OAI21X1_1817 ( .gnd(gnd), .vdd(vdd), .A(_1436_), .B(raddr2_0_bF_buf61_), .C(_4682_), .Y(_4683_) );
MUX2X1 MUX2X1_428 ( .gnd(gnd), .vdd(vdd), .A(_4683_), .B(_4681_), .S(raddr2_1_bF_buf9_), .Y(_4684_) );
NAND2X1 NAND2X1_866 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf4), .B(_4684_), .Y(_4685_) );
NAND2X1 NAND2X1_867 ( .gnd(gnd), .vdd(vdd), .A(regs_18__14_), .B(raddr2_0_bF_buf60_), .Y(_4686_) );
OAI21X1 OAI21X1_1818 ( .gnd(gnd), .vdd(vdd), .A(_1535_), .B(raddr2_0_bF_buf59_), .C(_4686_), .Y(_4687_) );
NAND2X1 NAND2X1_868 ( .gnd(gnd), .vdd(vdd), .A(regs_16__14_), .B(raddr2_0_bF_buf58_), .Y(_4688_) );
OAI21X1 OAI21X1_1819 ( .gnd(gnd), .vdd(vdd), .A(_1633_), .B(raddr2_0_bF_buf57_), .C(_4688_), .Y(_4689_) );
MUX2X1 MUX2X1_429 ( .gnd(gnd), .vdd(vdd), .A(_4689_), .B(_4687_), .S(raddr2_1_bF_buf8_), .Y(_4690_) );
AOI21X1 AOI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(raddr2_2_bF_buf0_), .B(_4690_), .C(_4033__bF_buf7), .Y(_4691_) );
OAI21X1 OAI21X1_1820 ( .gnd(gnd), .vdd(vdd), .A(_1171_), .B(raddr2_0_bF_buf56_), .C(raddr2_2_bF_buf10_), .Y(_4692_) );
AOI21X1 AOI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(regs_26__14_), .B(raddr2_0_bF_buf55_), .C(_4692_), .Y(_4693_) );
OAI21X1 OAI21X1_1821 ( .gnd(gnd), .vdd(vdd), .A(regs_30__14_), .B(raddr2_2_bF_buf9_), .C(_4038__bF_buf8), .Y(_4694_) );
OAI21X1 OAI21X1_1822 ( .gnd(gnd), .vdd(vdd), .A(_3130_), .B(raddr2_0_bF_buf54_), .C(raddr2_2_bF_buf8_), .Y(_4695_) );
AOI21X1 AOI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(regs_24__14_), .B(raddr2_0_bF_buf53_), .C(_4695_), .Y(_4696_) );
NOR2X1 NOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf52_), .B(_3133_), .Y(_4697_) );
NAND2X1 NAND2X1_869 ( .gnd(gnd), .vdd(vdd), .A(regs_28__14_), .B(raddr2_0_bF_buf51_), .Y(_4698_) );
NAND2X1 NAND2X1_870 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf3), .B(_4698_), .Y(_4699_) );
OAI21X1 OAI21X1_1823 ( .gnd(gnd), .vdd(vdd), .A(_4699_), .B(_4697_), .C(raddr2_1_bF_buf7_), .Y(_4700_) );
OAI22X1 OAI22X1_78 ( .gnd(gnd), .vdd(vdd), .A(_4693_), .B(_4694_), .C(_4700_), .D(_4696_), .Y(_4701_) );
AOI22X1 AOI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_4701_), .B(_4033__bF_buf6), .C(_4685_), .D(_4691_), .Y(_4702_) );
OAI21X1 OAI21X1_1824 ( .gnd(gnd), .vdd(vdd), .A(_3140_), .B(raddr2_0_bF_buf50_), .C(raddr2_1_bF_buf6_), .Y(_4703_) );
AOI21X1 AOI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(regs_4__14_), .B(raddr2_0_bF_buf49_), .C(_4703_), .Y(_4704_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(regs_6__14_), .B(raddr2_0_bF_buf48_), .Y(_4705_) );
OAI21X1 OAI21X1_1825 ( .gnd(gnd), .vdd(vdd), .A(_2129_), .B(raddr2_0_bF_buf47_), .C(_4038__bF_buf7), .Y(_4706_) );
OAI21X1 OAI21X1_1826 ( .gnd(gnd), .vdd(vdd), .A(_4706_), .B(_4705_), .C(_4036__bF_buf2), .Y(_4707_) );
OAI21X1 OAI21X1_1827 ( .gnd(gnd), .vdd(vdd), .A(_3146_), .B(raddr2_0_bF_buf46_), .C(raddr2_1_bF_buf5_), .Y(_4708_) );
AOI21X1 AOI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(regs_0__14_), .B(raddr2_0_bF_buf45_), .C(_4708_), .Y(_4709_) );
NOR2X1 NOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf44_), .B(_3149_), .Y(_4710_) );
NAND2X1 NAND2X1_871 ( .gnd(gnd), .vdd(vdd), .A(regs_2__14_), .B(raddr2_0_bF_buf43_), .Y(_4711_) );
NAND2X1 NAND2X1_872 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf6), .B(_4711_), .Y(_4712_) );
OAI21X1 OAI21X1_1828 ( .gnd(gnd), .vdd(vdd), .A(_4712_), .B(_4710_), .C(raddr2_2_bF_buf7_), .Y(_4713_) );
OAI22X1 OAI22X1_79 ( .gnd(gnd), .vdd(vdd), .A(_4709_), .B(_4713_), .C(_4707_), .D(_4704_), .Y(_4714_) );
NAND2X1 NAND2X1_873 ( .gnd(gnd), .vdd(vdd), .A(regs_10__14_), .B(raddr2_0_bF_buf42_), .Y(_4715_) );
OAI21X1 OAI21X1_1829 ( .gnd(gnd), .vdd(vdd), .A(_1930_), .B(raddr2_0_bF_buf41_), .C(_4715_), .Y(_4716_) );
NAND2X1 NAND2X1_874 ( .gnd(gnd), .vdd(vdd), .A(regs_8__14_), .B(raddr2_0_bF_buf40_), .Y(_4717_) );
OAI21X1 OAI21X1_1830 ( .gnd(gnd), .vdd(vdd), .A(_2028_), .B(raddr2_0_bF_buf39_), .C(_4717_), .Y(_4718_) );
MUX2X1 MUX2X1_430 ( .gnd(gnd), .vdd(vdd), .A(_4718_), .B(_4716_), .S(raddr2_1_bF_buf4_), .Y(_4719_) );
NAND2X1 NAND2X1_875 ( .gnd(gnd), .vdd(vdd), .A(regs_14__14_), .B(raddr2_0_bF_buf38_), .Y(_4720_) );
OAI21X1 OAI21X1_1831 ( .gnd(gnd), .vdd(vdd), .A(_1733_), .B(raddr2_0_bF_buf37_), .C(_4720_), .Y(_4721_) );
NAND2X1 NAND2X1_876 ( .gnd(gnd), .vdd(vdd), .A(regs_12__14_), .B(raddr2_0_bF_buf36_), .Y(_4722_) );
OAI21X1 OAI21X1_1832 ( .gnd(gnd), .vdd(vdd), .A(_1831_), .B(raddr2_0_bF_buf35_), .C(_4722_), .Y(_4723_) );
MUX2X1 MUX2X1_431 ( .gnd(gnd), .vdd(vdd), .A(_4723_), .B(_4721_), .S(raddr2_1_bF_buf3_), .Y(_4724_) );
MUX2X1 MUX2X1_432 ( .gnd(gnd), .vdd(vdd), .A(_4724_), .B(_4719_), .S(_4036__bF_buf1), .Y(_4725_) );
MUX2X1 MUX2X1_433 ( .gnd(gnd), .vdd(vdd), .A(_4725_), .B(_4714_), .S(_4033__bF_buf5), .Y(_4726_) );
MUX2X1 MUX2X1_434 ( .gnd(gnd), .vdd(vdd), .A(_4726_), .B(_4702_), .S(raddr2_4_bF_buf0_), .Y(_5512__14_) );
NAND2X1 NAND2X1_877 ( .gnd(gnd), .vdd(vdd), .A(regs_22__15_), .B(raddr2_0_bF_buf34_), .Y(_4727_) );
OAI21X1 OAI21X1_1833 ( .gnd(gnd), .vdd(vdd), .A(_1340_), .B(raddr2_0_bF_buf33_), .C(_4727_), .Y(_4728_) );
NAND2X1 NAND2X1_878 ( .gnd(gnd), .vdd(vdd), .A(regs_20__15_), .B(raddr2_0_bF_buf32_), .Y(_4729_) );
OAI21X1 OAI21X1_1834 ( .gnd(gnd), .vdd(vdd), .A(_1438_), .B(raddr2_0_bF_buf31_), .C(_4729_), .Y(_4730_) );
MUX2X1 MUX2X1_435 ( .gnd(gnd), .vdd(vdd), .A(_4730_), .B(_4728_), .S(raddr2_1_bF_buf2_), .Y(_4731_) );
NAND2X1 NAND2X1_879 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf0), .B(_4731_), .Y(_4732_) );
NAND2X1 NAND2X1_880 ( .gnd(gnd), .vdd(vdd), .A(regs_18__15_), .B(raddr2_0_bF_buf30_), .Y(_4733_) );
OAI21X1 OAI21X1_1835 ( .gnd(gnd), .vdd(vdd), .A(_1537_), .B(raddr2_0_bF_buf29_), .C(_4733_), .Y(_4734_) );
NAND2X1 NAND2X1_881 ( .gnd(gnd), .vdd(vdd), .A(regs_16__15_), .B(raddr2_0_bF_buf28_), .Y(_4735_) );
OAI21X1 OAI21X1_1836 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .B(raddr2_0_bF_buf27_), .C(_4735_), .Y(_4736_) );
MUX2X1 MUX2X1_436 ( .gnd(gnd), .vdd(vdd), .A(_4736_), .B(_4734_), .S(raddr2_1_bF_buf1_), .Y(_4737_) );
AOI21X1 AOI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(raddr2_2_bF_buf6_), .B(_4737_), .C(_4033__bF_buf4), .Y(_4738_) );
OAI21X1 OAI21X1_1837 ( .gnd(gnd), .vdd(vdd), .A(_1173_), .B(raddr2_0_bF_buf26_), .C(raddr2_2_bF_buf5_), .Y(_4739_) );
AOI21X1 AOI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(regs_26__15_), .B(raddr2_0_bF_buf25_), .C(_4739_), .Y(_4740_) );
OAI21X1 OAI21X1_1838 ( .gnd(gnd), .vdd(vdd), .A(regs_30__15_), .B(raddr2_2_bF_buf4_), .C(_4038__bF_buf5), .Y(_4741_) );
OAI21X1 OAI21X1_1839 ( .gnd(gnd), .vdd(vdd), .A(_3185_), .B(raddr2_0_bF_buf24_), .C(raddr2_2_bF_buf3_), .Y(_4742_) );
AOI21X1 AOI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(regs_24__15_), .B(raddr2_0_bF_buf23_), .C(_4742_), .Y(_4743_) );
NOR2X1 NOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf22_), .B(_3179_), .Y(_4744_) );
NAND2X1 NAND2X1_882 ( .gnd(gnd), .vdd(vdd), .A(regs_28__15_), .B(raddr2_0_bF_buf21_), .Y(_4745_) );
NAND2X1 NAND2X1_883 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf8), .B(_4745_), .Y(_4746_) );
OAI21X1 OAI21X1_1840 ( .gnd(gnd), .vdd(vdd), .A(_4746_), .B(_4744_), .C(raddr2_1_bF_buf0_), .Y(_4747_) );
OAI22X1 OAI22X1_80 ( .gnd(gnd), .vdd(vdd), .A(_4740_), .B(_4741_), .C(_4747_), .D(_4743_), .Y(_4748_) );
AOI22X1 AOI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_4748_), .B(_4033__bF_buf3), .C(_4732_), .D(_4738_), .Y(_4749_) );
OAI21X1 OAI21X1_1841 ( .gnd(gnd), .vdd(vdd), .A(_3193_), .B(raddr2_0_bF_buf20_), .C(raddr2_1_bF_buf14_bF_buf3_), .Y(_4750_) );
AOI21X1 AOI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(regs_4__15_), .B(raddr2_0_bF_buf19_), .C(_4750_), .Y(_4751_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(regs_6__15_), .B(raddr2_0_bF_buf18_), .Y(_4752_) );
OAI21X1 OAI21X1_1842 ( .gnd(gnd), .vdd(vdd), .A(_2131_), .B(raddr2_0_bF_buf17_), .C(_4038__bF_buf4), .Y(_4753_) );
OAI21X1 OAI21X1_1843 ( .gnd(gnd), .vdd(vdd), .A(_4753_), .B(_4752_), .C(_4036__bF_buf7), .Y(_4754_) );
OAI21X1 OAI21X1_1844 ( .gnd(gnd), .vdd(vdd), .A(_3200_), .B(raddr2_0_bF_buf16_), .C(raddr2_1_bF_buf13_bF_buf3_), .Y(_4755_) );
AOI21X1 AOI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(regs_0__15_), .B(raddr2_0_bF_buf15_), .C(_4755_), .Y(_4756_) );
NOR2X1 NOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf14_), .B(_3197_), .Y(_4757_) );
NAND2X1 NAND2X1_884 ( .gnd(gnd), .vdd(vdd), .A(regs_2__15_), .B(raddr2_0_bF_buf13_), .Y(_4758_) );
NAND2X1 NAND2X1_885 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf3), .B(_4758_), .Y(_4759_) );
OAI21X1 OAI21X1_1845 ( .gnd(gnd), .vdd(vdd), .A(_4759_), .B(_4757_), .C(raddr2_2_bF_buf2_), .Y(_4760_) );
OAI22X1 OAI22X1_81 ( .gnd(gnd), .vdd(vdd), .A(_4756_), .B(_4760_), .C(_4754_), .D(_4751_), .Y(_4761_) );
NAND2X1 NAND2X1_886 ( .gnd(gnd), .vdd(vdd), .A(regs_10__15_), .B(raddr2_0_bF_buf12_), .Y(_4762_) );
OAI21X1 OAI21X1_1846 ( .gnd(gnd), .vdd(vdd), .A(_1932_), .B(raddr2_0_bF_buf11_), .C(_4762_), .Y(_4763_) );
NAND2X1 NAND2X1_887 ( .gnd(gnd), .vdd(vdd), .A(regs_8__15_), .B(raddr2_0_bF_buf10_), .Y(_4764_) );
OAI21X1 OAI21X1_1847 ( .gnd(gnd), .vdd(vdd), .A(_2030_), .B(raddr2_0_bF_buf9_), .C(_4764_), .Y(_4765_) );
MUX2X1 MUX2X1_437 ( .gnd(gnd), .vdd(vdd), .A(_4765_), .B(_4763_), .S(raddr2_1_bF_buf12_bF_buf3_), .Y(_4766_) );
NAND2X1 NAND2X1_888 ( .gnd(gnd), .vdd(vdd), .A(regs_14__15_), .B(raddr2_0_bF_buf8_), .Y(_4767_) );
OAI21X1 OAI21X1_1848 ( .gnd(gnd), .vdd(vdd), .A(_1735_), .B(raddr2_0_bF_buf7_), .C(_4767_), .Y(_4768_) );
NAND2X1 NAND2X1_889 ( .gnd(gnd), .vdd(vdd), .A(regs_12__15_), .B(raddr2_0_bF_buf6_), .Y(_4769_) );
OAI21X1 OAI21X1_1849 ( .gnd(gnd), .vdd(vdd), .A(_1833_), .B(raddr2_0_bF_buf5_), .C(_4769_), .Y(_4770_) );
MUX2X1 MUX2X1_438 ( .gnd(gnd), .vdd(vdd), .A(_4770_), .B(_4768_), .S(raddr2_1_bF_buf11_), .Y(_4771_) );
MUX2X1 MUX2X1_439 ( .gnd(gnd), .vdd(vdd), .A(_4771_), .B(_4766_), .S(_4036__bF_buf6), .Y(_4772_) );
MUX2X1 MUX2X1_440 ( .gnd(gnd), .vdd(vdd), .A(_4772_), .B(_4761_), .S(_4033__bF_buf2), .Y(_4773_) );
MUX2X1 MUX2X1_441 ( .gnd(gnd), .vdd(vdd), .A(_4773_), .B(_4749_), .S(raddr2_4_bF_buf4_), .Y(_5512__15_) );
NAND2X1 NAND2X1_890 ( .gnd(gnd), .vdd(vdd), .A(regs_22__16_), .B(raddr2_0_bF_buf4_), .Y(_4774_) );
OAI21X1 OAI21X1_1850 ( .gnd(gnd), .vdd(vdd), .A(_1342_), .B(raddr2_0_bF_buf3_), .C(_4774_), .Y(_4775_) );
NAND2X1 NAND2X1_891 ( .gnd(gnd), .vdd(vdd), .A(regs_20__16_), .B(raddr2_0_bF_buf2_), .Y(_4776_) );
OAI21X1 OAI21X1_1851 ( .gnd(gnd), .vdd(vdd), .A(_1440_), .B(raddr2_0_bF_buf1_), .C(_4776_), .Y(_4777_) );
MUX2X1 MUX2X1_442 ( .gnd(gnd), .vdd(vdd), .A(_4777_), .B(_4775_), .S(raddr2_1_bF_buf10_), .Y(_4778_) );
NAND2X1 NAND2X1_892 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf5), .B(_4778_), .Y(_4779_) );
NAND2X1 NAND2X1_893 ( .gnd(gnd), .vdd(vdd), .A(regs_18__16_), .B(raddr2_0_bF_buf0_), .Y(_4780_) );
OAI21X1 OAI21X1_1852 ( .gnd(gnd), .vdd(vdd), .A(_1539_), .B(raddr2_0_bF_buf96_), .C(_4780_), .Y(_4781_) );
NAND2X1 NAND2X1_894 ( .gnd(gnd), .vdd(vdd), .A(regs_16__16_), .B(raddr2_0_bF_buf95_), .Y(_4782_) );
OAI21X1 OAI21X1_1853 ( .gnd(gnd), .vdd(vdd), .A(_1637_), .B(raddr2_0_bF_buf94_), .C(_4782_), .Y(_4783_) );
MUX2X1 MUX2X1_443 ( .gnd(gnd), .vdd(vdd), .A(_4783_), .B(_4781_), .S(raddr2_1_bF_buf9_), .Y(_4784_) );
AOI21X1 AOI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(raddr2_2_bF_buf1_), .B(_4784_), .C(_4033__bF_buf1), .Y(_4785_) );
OAI21X1 OAI21X1_1854 ( .gnd(gnd), .vdd(vdd), .A(_1175_), .B(raddr2_0_bF_buf93_), .C(raddr2_2_bF_buf0_), .Y(_4786_) );
AOI21X1 AOI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(regs_26__16_), .B(raddr2_0_bF_buf92_), .C(_4786_), .Y(_4787_) );
OAI21X1 OAI21X1_1855 ( .gnd(gnd), .vdd(vdd), .A(regs_30__16_), .B(raddr2_2_bF_buf10_), .C(_4038__bF_buf2), .Y(_4788_) );
OAI21X1 OAI21X1_1856 ( .gnd(gnd), .vdd(vdd), .A(_3232_), .B(raddr2_0_bF_buf91_), .C(raddr2_2_bF_buf9_), .Y(_4789_) );
AOI21X1 AOI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(regs_24__16_), .B(raddr2_0_bF_buf90_), .C(_4789_), .Y(_4790_) );
NOR2X1 NOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf89_), .B(_3235_), .Y(_4791_) );
NAND2X1 NAND2X1_895 ( .gnd(gnd), .vdd(vdd), .A(regs_28__16_), .B(raddr2_0_bF_buf88_), .Y(_4792_) );
NAND2X1 NAND2X1_896 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf4), .B(_4792_), .Y(_4793_) );
OAI21X1 OAI21X1_1857 ( .gnd(gnd), .vdd(vdd), .A(_4793_), .B(_4791_), .C(raddr2_1_bF_buf8_), .Y(_4794_) );
OAI22X1 OAI22X1_82 ( .gnd(gnd), .vdd(vdd), .A(_4787_), .B(_4788_), .C(_4794_), .D(_4790_), .Y(_4795_) );
AOI22X1 AOI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_4795_), .B(_4033__bF_buf0), .C(_4779_), .D(_4785_), .Y(_4796_) );
OAI21X1 OAI21X1_1858 ( .gnd(gnd), .vdd(vdd), .A(_3242_), .B(raddr2_0_bF_buf87_), .C(raddr2_1_bF_buf7_), .Y(_4797_) );
AOI21X1 AOI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(regs_4__16_), .B(raddr2_0_bF_buf86_), .C(_4797_), .Y(_4798_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(regs_6__16_), .B(raddr2_0_bF_buf85_), .Y(_4799_) );
OAI21X1 OAI21X1_1859 ( .gnd(gnd), .vdd(vdd), .A(_2133_), .B(raddr2_0_bF_buf84_), .C(_4038__bF_buf1), .Y(_4800_) );
OAI21X1 OAI21X1_1860 ( .gnd(gnd), .vdd(vdd), .A(_4800_), .B(_4799_), .C(_4036__bF_buf3), .Y(_4801_) );
OAI21X1 OAI21X1_1861 ( .gnd(gnd), .vdd(vdd), .A(_3248_), .B(raddr2_0_bF_buf83_), .C(raddr2_1_bF_buf6_), .Y(_4802_) );
AOI21X1 AOI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(regs_0__16_), .B(raddr2_0_bF_buf82_), .C(_4802_), .Y(_4803_) );
NOR2X1 NOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf81_), .B(_3251_), .Y(_4804_) );
NAND2X1 NAND2X1_897 ( .gnd(gnd), .vdd(vdd), .A(regs_2__16_), .B(raddr2_0_bF_buf80_), .Y(_4805_) );
NAND2X1 NAND2X1_898 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf0), .B(_4805_), .Y(_4806_) );
OAI21X1 OAI21X1_1862 ( .gnd(gnd), .vdd(vdd), .A(_4806_), .B(_4804_), .C(raddr2_2_bF_buf8_), .Y(_4807_) );
OAI22X1 OAI22X1_83 ( .gnd(gnd), .vdd(vdd), .A(_4803_), .B(_4807_), .C(_4801_), .D(_4798_), .Y(_4808_) );
NAND2X1 NAND2X1_899 ( .gnd(gnd), .vdd(vdd), .A(regs_10__16_), .B(raddr2_0_bF_buf79_), .Y(_4809_) );
OAI21X1 OAI21X1_1863 ( .gnd(gnd), .vdd(vdd), .A(_1934_), .B(raddr2_0_bF_buf78_), .C(_4809_), .Y(_4810_) );
NAND2X1 NAND2X1_900 ( .gnd(gnd), .vdd(vdd), .A(regs_8__16_), .B(raddr2_0_bF_buf77_), .Y(_4811_) );
OAI21X1 OAI21X1_1864 ( .gnd(gnd), .vdd(vdd), .A(_2032_), .B(raddr2_0_bF_buf76_), .C(_4811_), .Y(_4812_) );
MUX2X1 MUX2X1_444 ( .gnd(gnd), .vdd(vdd), .A(_4812_), .B(_4810_), .S(raddr2_1_bF_buf5_), .Y(_4813_) );
NAND2X1 NAND2X1_901 ( .gnd(gnd), .vdd(vdd), .A(regs_14__16_), .B(raddr2_0_bF_buf75_), .Y(_4814_) );
OAI21X1 OAI21X1_1865 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(raddr2_0_bF_buf74_), .C(_4814_), .Y(_4815_) );
NAND2X1 NAND2X1_902 ( .gnd(gnd), .vdd(vdd), .A(regs_12__16_), .B(raddr2_0_bF_buf73_), .Y(_4816_) );
OAI21X1 OAI21X1_1866 ( .gnd(gnd), .vdd(vdd), .A(_1835_), .B(raddr2_0_bF_buf72_), .C(_4816_), .Y(_4817_) );
MUX2X1 MUX2X1_445 ( .gnd(gnd), .vdd(vdd), .A(_4817_), .B(_4815_), .S(raddr2_1_bF_buf4_), .Y(_4818_) );
MUX2X1 MUX2X1_446 ( .gnd(gnd), .vdd(vdd), .A(_4818_), .B(_4813_), .S(_4036__bF_buf2), .Y(_4819_) );
MUX2X1 MUX2X1_447 ( .gnd(gnd), .vdd(vdd), .A(_4819_), .B(_4808_), .S(_4033__bF_buf7), .Y(_4820_) );
MUX2X1 MUX2X1_448 ( .gnd(gnd), .vdd(vdd), .A(_4820_), .B(_4796_), .S(raddr2_4_bF_buf3_), .Y(_5512__16_) );
OAI21X1 OAI21X1_1867 ( .gnd(gnd), .vdd(vdd), .A(_1442_), .B(raddr2_0_bF_buf71_), .C(raddr2_1_bF_buf3_), .Y(_4821_) );
AOI21X1 AOI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(regs_20__17_), .B(raddr2_0_bF_buf70_), .C(_4821_), .Y(_4822_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(regs_22__17_), .B(raddr2_0_bF_buf69_), .Y(_4823_) );
OAI21X1 OAI21X1_1868 ( .gnd(gnd), .vdd(vdd), .A(_1344_), .B(raddr2_0_bF_buf68_), .C(_4038__bF_buf8), .Y(_4824_) );
OAI21X1 OAI21X1_1869 ( .gnd(gnd), .vdd(vdd), .A(_4824_), .B(_4823_), .C(_4036__bF_buf1), .Y(_4825_) );
OAI21X1 OAI21X1_1870 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .B(raddr2_0_bF_buf67_), .C(raddr2_1_bF_buf2_), .Y(_4826_) );
AOI21X1 AOI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(regs_16__17_), .B(raddr2_0_bF_buf66_), .C(_4826_), .Y(_4827_) );
NOR2X1 NOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf65_), .B(_1541_), .Y(_4828_) );
NAND2X1 NAND2X1_903 ( .gnd(gnd), .vdd(vdd), .A(regs_18__17_), .B(raddr2_0_bF_buf64_), .Y(_4829_) );
NAND2X1 NAND2X1_904 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf7), .B(_4829_), .Y(_4830_) );
OAI21X1 OAI21X1_1871 ( .gnd(gnd), .vdd(vdd), .A(_4830_), .B(_4828_), .C(raddr2_2_bF_buf7_), .Y(_4831_) );
OAI22X1 OAI22X1_84 ( .gnd(gnd), .vdd(vdd), .A(_4827_), .B(_4831_), .C(_4825_), .D(_4822_), .Y(_4832_) );
NAND2X1 NAND2X1_905 ( .gnd(gnd), .vdd(vdd), .A(regs_28__17_), .B(raddr2_0_bF_buf63_), .Y(_4833_) );
OAI21X1 OAI21X1_1872 ( .gnd(gnd), .vdd(vdd), .A(_3287_), .B(raddr2_0_bF_buf62_), .C(_4833_), .Y(_4834_) );
MUX2X1 MUX2X1_449 ( .gnd(gnd), .vdd(vdd), .A(_4834_), .B(regs_30__17_), .S(raddr2_1_bF_buf1_), .Y(_4835_) );
NAND2X1 NAND2X1_906 ( .gnd(gnd), .vdd(vdd), .A(regs_26__17_), .B(raddr2_0_bF_buf61_), .Y(_4836_) );
OAI21X1 OAI21X1_1873 ( .gnd(gnd), .vdd(vdd), .A(_1177_), .B(raddr2_0_bF_buf60_), .C(_4836_), .Y(_4837_) );
NAND2X1 NAND2X1_907 ( .gnd(gnd), .vdd(vdd), .A(regs_24__17_), .B(raddr2_0_bF_buf59_), .Y(_4838_) );
OAI21X1 OAI21X1_1874 ( .gnd(gnd), .vdd(vdd), .A(_3284_), .B(raddr2_0_bF_buf58_), .C(_4838_), .Y(_4839_) );
MUX2X1 MUX2X1_450 ( .gnd(gnd), .vdd(vdd), .A(_4839_), .B(_4837_), .S(raddr2_1_bF_buf0_), .Y(_4840_) );
MUX2X1 MUX2X1_451 ( .gnd(gnd), .vdd(vdd), .A(_4840_), .B(_4835_), .S(raddr2_2_bF_buf6_), .Y(_4841_) );
MUX2X1 MUX2X1_452 ( .gnd(gnd), .vdd(vdd), .A(_4841_), .B(_4832_), .S(_4033__bF_buf6), .Y(_4842_) );
NAND2X1 NAND2X1_908 ( .gnd(gnd), .vdd(vdd), .A(regs_6__17_), .B(raddr2_0_bF_buf57_), .Y(_4843_) );
OAI21X1 OAI21X1_1875 ( .gnd(gnd), .vdd(vdd), .A(_2135_), .B(raddr2_0_bF_buf56_), .C(_4843_), .Y(_4844_) );
NAND2X1 NAND2X1_909 ( .gnd(gnd), .vdd(vdd), .A(regs_4__17_), .B(raddr2_0_bF_buf55_), .Y(_4845_) );
OAI21X1 OAI21X1_1876 ( .gnd(gnd), .vdd(vdd), .A(_3294_), .B(raddr2_0_bF_buf54_), .C(_4845_), .Y(_4846_) );
MUX2X1 MUX2X1_453 ( .gnd(gnd), .vdd(vdd), .A(_4846_), .B(_4844_), .S(raddr2_1_bF_buf14_bF_buf2_), .Y(_4847_) );
NAND2X1 NAND2X1_910 ( .gnd(gnd), .vdd(vdd), .A(regs_2__17_), .B(raddr2_0_bF_buf53_), .Y(_4848_) );
OAI21X1 OAI21X1_1877 ( .gnd(gnd), .vdd(vdd), .A(_3303_), .B(raddr2_0_bF_buf52_), .C(_4848_), .Y(_4849_) );
NAND2X1 NAND2X1_911 ( .gnd(gnd), .vdd(vdd), .A(regs_0__17_), .B(raddr2_0_bF_buf51_), .Y(_4850_) );
OAI21X1 OAI21X1_1878 ( .gnd(gnd), .vdd(vdd), .A(_3300_), .B(raddr2_0_bF_buf50_), .C(_4850_), .Y(_4851_) );
MUX2X1 MUX2X1_454 ( .gnd(gnd), .vdd(vdd), .A(_4851_), .B(_4849_), .S(raddr2_1_bF_buf13_bF_buf2_), .Y(_4852_) );
MUX2X1 MUX2X1_455 ( .gnd(gnd), .vdd(vdd), .A(_4852_), .B(_4847_), .S(raddr2_2_bF_buf5_), .Y(_4853_) );
NAND2X1 NAND2X1_912 ( .gnd(gnd), .vdd(vdd), .A(regs_14__17_), .B(raddr2_0_bF_buf49_), .Y(_4854_) );
OAI21X1 OAI21X1_1879 ( .gnd(gnd), .vdd(vdd), .A(_1739_), .B(raddr2_0_bF_buf48_), .C(_4854_), .Y(_4855_) );
NAND2X1 NAND2X1_913 ( .gnd(gnd), .vdd(vdd), .A(regs_12__17_), .B(raddr2_0_bF_buf47_), .Y(_4856_) );
OAI21X1 OAI21X1_1880 ( .gnd(gnd), .vdd(vdd), .A(_1837_), .B(raddr2_0_bF_buf46_), .C(_4856_), .Y(_4857_) );
MUX2X1 MUX2X1_456 ( .gnd(gnd), .vdd(vdd), .A(_4857_), .B(_4855_), .S(raddr2_1_bF_buf12_bF_buf2_), .Y(_4858_) );
NAND2X1 NAND2X1_914 ( .gnd(gnd), .vdd(vdd), .A(regs_10__17_), .B(raddr2_0_bF_buf45_), .Y(_4859_) );
OAI21X1 OAI21X1_1881 ( .gnd(gnd), .vdd(vdd), .A(_1936_), .B(raddr2_0_bF_buf44_), .C(_4859_), .Y(_4860_) );
NAND2X1 NAND2X1_915 ( .gnd(gnd), .vdd(vdd), .A(regs_8__17_), .B(raddr2_0_bF_buf43_), .Y(_4861_) );
OAI21X1 OAI21X1_1882 ( .gnd(gnd), .vdd(vdd), .A(_2034_), .B(raddr2_0_bF_buf42_), .C(_4861_), .Y(_4862_) );
MUX2X1 MUX2X1_457 ( .gnd(gnd), .vdd(vdd), .A(_4862_), .B(_4860_), .S(raddr2_1_bF_buf11_), .Y(_4863_) );
MUX2X1 MUX2X1_458 ( .gnd(gnd), .vdd(vdd), .A(_4863_), .B(_4858_), .S(raddr2_2_bF_buf4_), .Y(_4864_) );
MUX2X1 MUX2X1_459 ( .gnd(gnd), .vdd(vdd), .A(_4864_), .B(_4853_), .S(_4033__bF_buf5), .Y(_4865_) );
MUX2X1 MUX2X1_460 ( .gnd(gnd), .vdd(vdd), .A(_4865_), .B(_4842_), .S(raddr2_4_bF_buf2_), .Y(_5512__17_) );
NAND2X1 NAND2X1_916 ( .gnd(gnd), .vdd(vdd), .A(regs_22__18_), .B(raddr2_0_bF_buf41_), .Y(_4866_) );
OAI21X1 OAI21X1_1883 ( .gnd(gnd), .vdd(vdd), .A(_1346_), .B(raddr2_0_bF_buf40_), .C(_4866_), .Y(_4867_) );
NAND2X1 NAND2X1_917 ( .gnd(gnd), .vdd(vdd), .A(regs_20__18_), .B(raddr2_0_bF_buf39_), .Y(_4868_) );
OAI21X1 OAI21X1_1884 ( .gnd(gnd), .vdd(vdd), .A(_1444_), .B(raddr2_0_bF_buf38_), .C(_4868_), .Y(_4869_) );
MUX2X1 MUX2X1_461 ( .gnd(gnd), .vdd(vdd), .A(_4869_), .B(_4867_), .S(raddr2_1_bF_buf10_), .Y(_4870_) );
NAND2X1 NAND2X1_918 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf0), .B(_4870_), .Y(_4871_) );
NAND2X1 NAND2X1_919 ( .gnd(gnd), .vdd(vdd), .A(regs_18__18_), .B(raddr2_0_bF_buf37_), .Y(_4872_) );
OAI21X1 OAI21X1_1885 ( .gnd(gnd), .vdd(vdd), .A(_1543_), .B(raddr2_0_bF_buf36_), .C(_4872_), .Y(_4873_) );
NAND2X1 NAND2X1_920 ( .gnd(gnd), .vdd(vdd), .A(regs_16__18_), .B(raddr2_0_bF_buf35_), .Y(_4874_) );
OAI21X1 OAI21X1_1886 ( .gnd(gnd), .vdd(vdd), .A(_1641_), .B(raddr2_0_bF_buf34_), .C(_4874_), .Y(_4875_) );
MUX2X1 MUX2X1_462 ( .gnd(gnd), .vdd(vdd), .A(_4875_), .B(_4873_), .S(raddr2_1_bF_buf9_), .Y(_4876_) );
AOI21X1 AOI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(raddr2_2_bF_buf3_), .B(_4876_), .C(_4033__bF_buf4), .Y(_4877_) );
OAI21X1 OAI21X1_1887 ( .gnd(gnd), .vdd(vdd), .A(_1179_), .B(raddr2_0_bF_buf33_), .C(raddr2_2_bF_buf2_), .Y(_4878_) );
AOI21X1 AOI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(regs_26__18_), .B(raddr2_0_bF_buf32_), .C(_4878_), .Y(_4879_) );
OAI21X1 OAI21X1_1888 ( .gnd(gnd), .vdd(vdd), .A(regs_30__18_), .B(raddr2_2_bF_buf1_), .C(_4038__bF_buf6), .Y(_4880_) );
OAI21X1 OAI21X1_1889 ( .gnd(gnd), .vdd(vdd), .A(_3366_), .B(raddr2_0_bF_buf31_), .C(raddr2_2_bF_buf0_), .Y(_4881_) );
AOI21X1 AOI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(regs_24__18_), .B(raddr2_0_bF_buf30_), .C(_4881_), .Y(_4882_) );
NOR2X1 NOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf29_), .B(_3360_), .Y(_4883_) );
NAND2X1 NAND2X1_921 ( .gnd(gnd), .vdd(vdd), .A(regs_28__18_), .B(raddr2_0_bF_buf28_), .Y(_4884_) );
NAND2X1 NAND2X1_922 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf8), .B(_4884_), .Y(_4885_) );
OAI21X1 OAI21X1_1890 ( .gnd(gnd), .vdd(vdd), .A(_4885_), .B(_4883_), .C(raddr2_1_bF_buf8_), .Y(_4886_) );
OAI22X1 OAI22X1_85 ( .gnd(gnd), .vdd(vdd), .A(_4879_), .B(_4880_), .C(_4886_), .D(_4882_), .Y(_4887_) );
AOI22X1 AOI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_4887_), .B(_4033__bF_buf3), .C(_4871_), .D(_4877_), .Y(_4888_) );
NAND2X1 NAND2X1_923 ( .gnd(gnd), .vdd(vdd), .A(regs_6__18_), .B(raddr2_0_bF_buf27_), .Y(_4889_) );
OAI21X1 OAI21X1_1891 ( .gnd(gnd), .vdd(vdd), .A(_2137_), .B(raddr2_0_bF_buf26_), .C(_4889_), .Y(_4890_) );
NAND2X1 NAND2X1_924 ( .gnd(gnd), .vdd(vdd), .A(regs_4__18_), .B(raddr2_0_bF_buf25_), .Y(_4891_) );
OAI21X1 OAI21X1_1892 ( .gnd(gnd), .vdd(vdd), .A(_3321_), .B(raddr2_0_bF_buf24_), .C(_4891_), .Y(_4892_) );
MUX2X1 MUX2X1_463 ( .gnd(gnd), .vdd(vdd), .A(_4892_), .B(_4890_), .S(raddr2_1_bF_buf7_), .Y(_4893_) );
NAND2X1 NAND2X1_925 ( .gnd(gnd), .vdd(vdd), .A(regs_2__18_), .B(raddr2_0_bF_buf23_), .Y(_4894_) );
OAI21X1 OAI21X1_1893 ( .gnd(gnd), .vdd(vdd), .A(_3330_), .B(raddr2_0_bF_buf22_), .C(_4894_), .Y(_4895_) );
NAND2X1 NAND2X1_926 ( .gnd(gnd), .vdd(vdd), .A(regs_0__18_), .B(raddr2_0_bF_buf21_), .Y(_4896_) );
OAI21X1 OAI21X1_1894 ( .gnd(gnd), .vdd(vdd), .A(_3327_), .B(raddr2_0_bF_buf20_), .C(_4896_), .Y(_4897_) );
MUX2X1 MUX2X1_464 ( .gnd(gnd), .vdd(vdd), .A(_4897_), .B(_4895_), .S(raddr2_1_bF_buf6_), .Y(_4898_) );
MUX2X1 MUX2X1_465 ( .gnd(gnd), .vdd(vdd), .A(_4898_), .B(_4893_), .S(raddr2_2_bF_buf10_), .Y(_4899_) );
NAND2X1 NAND2X1_927 ( .gnd(gnd), .vdd(vdd), .A(regs_10__18_), .B(raddr2_0_bF_buf19_), .Y(_4900_) );
OAI21X1 OAI21X1_1895 ( .gnd(gnd), .vdd(vdd), .A(_1938_), .B(raddr2_0_bF_buf18_), .C(_4900_), .Y(_4901_) );
NAND2X1 NAND2X1_928 ( .gnd(gnd), .vdd(vdd), .A(regs_8__18_), .B(raddr2_0_bF_buf17_), .Y(_4902_) );
OAI21X1 OAI21X1_1896 ( .gnd(gnd), .vdd(vdd), .A(_2036_), .B(raddr2_0_bF_buf16_), .C(_4902_), .Y(_4903_) );
MUX2X1 MUX2X1_466 ( .gnd(gnd), .vdd(vdd), .A(_4903_), .B(_4901_), .S(raddr2_1_bF_buf5_), .Y(_4904_) );
NAND2X1 NAND2X1_929 ( .gnd(gnd), .vdd(vdd), .A(regs_14__18_), .B(raddr2_0_bF_buf15_), .Y(_4905_) );
OAI21X1 OAI21X1_1897 ( .gnd(gnd), .vdd(vdd), .A(_1741_), .B(raddr2_0_bF_buf14_), .C(_4905_), .Y(_4906_) );
NAND2X1 NAND2X1_930 ( .gnd(gnd), .vdd(vdd), .A(regs_12__18_), .B(raddr2_0_bF_buf13_), .Y(_4907_) );
OAI21X1 OAI21X1_1898 ( .gnd(gnd), .vdd(vdd), .A(_1839_), .B(raddr2_0_bF_buf12_), .C(_4907_), .Y(_4908_) );
MUX2X1 MUX2X1_467 ( .gnd(gnd), .vdd(vdd), .A(_4908_), .B(_4906_), .S(raddr2_1_bF_buf4_), .Y(_4909_) );
MUX2X1 MUX2X1_468 ( .gnd(gnd), .vdd(vdd), .A(_4909_), .B(_4904_), .S(_4036__bF_buf7), .Y(_4910_) );
MUX2X1 MUX2X1_469 ( .gnd(gnd), .vdd(vdd), .A(_4910_), .B(_4899_), .S(_4033__bF_buf2), .Y(_4911_) );
MUX2X1 MUX2X1_470 ( .gnd(gnd), .vdd(vdd), .A(_4911_), .B(_4888_), .S(raddr2_4_bF_buf1_), .Y(_5512__18_) );
NAND2X1 NAND2X1_931 ( .gnd(gnd), .vdd(vdd), .A(regs_22__19_), .B(raddr2_0_bF_buf11_), .Y(_4912_) );
OAI21X1 OAI21X1_1899 ( .gnd(gnd), .vdd(vdd), .A(_1348_), .B(raddr2_0_bF_buf10_), .C(_4912_), .Y(_4913_) );
NAND2X1 NAND2X1_932 ( .gnd(gnd), .vdd(vdd), .A(regs_20__19_), .B(raddr2_0_bF_buf9_), .Y(_4914_) );
OAI21X1 OAI21X1_1900 ( .gnd(gnd), .vdd(vdd), .A(_1446_), .B(raddr2_0_bF_buf8_), .C(_4914_), .Y(_4915_) );
MUX2X1 MUX2X1_471 ( .gnd(gnd), .vdd(vdd), .A(_4915_), .B(_4913_), .S(raddr2_1_bF_buf3_), .Y(_4916_) );
NAND2X1 NAND2X1_933 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf6), .B(_4916_), .Y(_4917_) );
NAND2X1 NAND2X1_934 ( .gnd(gnd), .vdd(vdd), .A(regs_18__19_), .B(raddr2_0_bF_buf7_), .Y(_4918_) );
OAI21X1 OAI21X1_1901 ( .gnd(gnd), .vdd(vdd), .A(_1545_), .B(raddr2_0_bF_buf6_), .C(_4918_), .Y(_4919_) );
NAND2X1 NAND2X1_935 ( .gnd(gnd), .vdd(vdd), .A(regs_16__19_), .B(raddr2_0_bF_buf5_), .Y(_4920_) );
OAI21X1 OAI21X1_1902 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .B(raddr2_0_bF_buf4_), .C(_4920_), .Y(_4921_) );
MUX2X1 MUX2X1_472 ( .gnd(gnd), .vdd(vdd), .A(_4921_), .B(_4919_), .S(raddr2_1_bF_buf2_), .Y(_4922_) );
AOI21X1 AOI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(raddr2_2_bF_buf9_), .B(_4922_), .C(_4033__bF_buf1), .Y(_4923_) );
OAI21X1 OAI21X1_1903 ( .gnd(gnd), .vdd(vdd), .A(_1181_), .B(raddr2_0_bF_buf3_), .C(raddr2_2_bF_buf8_), .Y(_4924_) );
AOI21X1 AOI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(regs_26__19_), .B(raddr2_0_bF_buf2_), .C(_4924_), .Y(_4925_) );
OAI21X1 OAI21X1_1904 ( .gnd(gnd), .vdd(vdd), .A(regs_30__19_), .B(raddr2_2_bF_buf7_), .C(_4038__bF_buf5), .Y(_4926_) );
OAI21X1 OAI21X1_1905 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .B(raddr2_0_bF_buf1_), .C(raddr2_2_bF_buf6_), .Y(_4927_) );
AOI21X1 AOI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(regs_24__19_), .B(raddr2_0_bF_buf0_), .C(_4927_), .Y(_4928_) );
NOR2X1 NOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf96_), .B(_3390_), .Y(_4929_) );
NAND2X1 NAND2X1_936 ( .gnd(gnd), .vdd(vdd), .A(regs_28__19_), .B(raddr2_0_bF_buf95_), .Y(_4930_) );
NAND2X1 NAND2X1_937 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf5), .B(_4930_), .Y(_4931_) );
OAI21X1 OAI21X1_1906 ( .gnd(gnd), .vdd(vdd), .A(_4931_), .B(_4929_), .C(raddr2_1_bF_buf1_), .Y(_4932_) );
OAI22X1 OAI22X1_86 ( .gnd(gnd), .vdd(vdd), .A(_4925_), .B(_4926_), .C(_4932_), .D(_4928_), .Y(_4933_) );
AOI22X1 AOI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_4933_), .B(_4033__bF_buf0), .C(_4917_), .D(_4923_), .Y(_4934_) );
NAND2X1 NAND2X1_938 ( .gnd(gnd), .vdd(vdd), .A(regs_6__19_), .B(raddr2_0_bF_buf94_), .Y(_4935_) );
OAI21X1 OAI21X1_1907 ( .gnd(gnd), .vdd(vdd), .A(_2139_), .B(raddr2_0_bF_buf93_), .C(_4935_), .Y(_4936_) );
NAND2X1 NAND2X1_939 ( .gnd(gnd), .vdd(vdd), .A(regs_4__19_), .B(raddr2_0_bF_buf92_), .Y(_4937_) );
OAI21X1 OAI21X1_1908 ( .gnd(gnd), .vdd(vdd), .A(_3399_), .B(raddr2_0_bF_buf91_), .C(_4937_), .Y(_4938_) );
MUX2X1 MUX2X1_473 ( .gnd(gnd), .vdd(vdd), .A(_4938_), .B(_4936_), .S(raddr2_1_bF_buf0_), .Y(_4939_) );
NAND2X1 NAND2X1_940 ( .gnd(gnd), .vdd(vdd), .A(regs_2__19_), .B(raddr2_0_bF_buf90_), .Y(_4940_) );
OAI21X1 OAI21X1_1909 ( .gnd(gnd), .vdd(vdd), .A(_3403_), .B(raddr2_0_bF_buf89_), .C(_4940_), .Y(_4941_) );
NAND2X1 NAND2X1_941 ( .gnd(gnd), .vdd(vdd), .A(regs_0__19_), .B(raddr2_0_bF_buf88_), .Y(_4942_) );
OAI21X1 OAI21X1_1910 ( .gnd(gnd), .vdd(vdd), .A(_3406_), .B(raddr2_0_bF_buf87_), .C(_4942_), .Y(_4943_) );
MUX2X1 MUX2X1_474 ( .gnd(gnd), .vdd(vdd), .A(_4943_), .B(_4941_), .S(raddr2_1_bF_buf14_bF_buf1_), .Y(_4944_) );
MUX2X1 MUX2X1_475 ( .gnd(gnd), .vdd(vdd), .A(_4944_), .B(_4939_), .S(raddr2_2_bF_buf5_), .Y(_4945_) );
NAND2X1 NAND2X1_942 ( .gnd(gnd), .vdd(vdd), .A(regs_10__19_), .B(raddr2_0_bF_buf86_), .Y(_4946_) );
OAI21X1 OAI21X1_1911 ( .gnd(gnd), .vdd(vdd), .A(_1940_), .B(raddr2_0_bF_buf85_), .C(_4946_), .Y(_4947_) );
NAND2X1 NAND2X1_943 ( .gnd(gnd), .vdd(vdd), .A(regs_8__19_), .B(raddr2_0_bF_buf84_), .Y(_4948_) );
OAI21X1 OAI21X1_1912 ( .gnd(gnd), .vdd(vdd), .A(_2038_), .B(raddr2_0_bF_buf83_), .C(_4948_), .Y(_4949_) );
MUX2X1 MUX2X1_476 ( .gnd(gnd), .vdd(vdd), .A(_4949_), .B(_4947_), .S(raddr2_1_bF_buf13_bF_buf1_), .Y(_4950_) );
NAND2X1 NAND2X1_944 ( .gnd(gnd), .vdd(vdd), .A(regs_14__19_), .B(raddr2_0_bF_buf82_), .Y(_4951_) );
OAI21X1 OAI21X1_1913 ( .gnd(gnd), .vdd(vdd), .A(_1743_), .B(raddr2_0_bF_buf81_), .C(_4951_), .Y(_4952_) );
NAND2X1 NAND2X1_945 ( .gnd(gnd), .vdd(vdd), .A(regs_12__19_), .B(raddr2_0_bF_buf80_), .Y(_4953_) );
OAI21X1 OAI21X1_1914 ( .gnd(gnd), .vdd(vdd), .A(_1841_), .B(raddr2_0_bF_buf79_), .C(_4953_), .Y(_4954_) );
MUX2X1 MUX2X1_477 ( .gnd(gnd), .vdd(vdd), .A(_4954_), .B(_4952_), .S(raddr2_1_bF_buf12_bF_buf1_), .Y(_4955_) );
MUX2X1 MUX2X1_478 ( .gnd(gnd), .vdd(vdd), .A(_4955_), .B(_4950_), .S(_4036__bF_buf4), .Y(_4956_) );
MUX2X1 MUX2X1_479 ( .gnd(gnd), .vdd(vdd), .A(_4956_), .B(_4945_), .S(_4033__bF_buf7), .Y(_4957_) );
MUX2X1 MUX2X1_480 ( .gnd(gnd), .vdd(vdd), .A(_4957_), .B(_4934_), .S(raddr2_4_bF_buf0_), .Y(_5512__19_) );
NAND2X1 NAND2X1_946 ( .gnd(gnd), .vdd(vdd), .A(regs_22__20_), .B(raddr2_0_bF_buf78_), .Y(_4958_) );
OAI21X1 OAI21X1_1915 ( .gnd(gnd), .vdd(vdd), .A(_1350_), .B(raddr2_0_bF_buf77_), .C(_4958_), .Y(_4959_) );
NAND2X1 NAND2X1_947 ( .gnd(gnd), .vdd(vdd), .A(regs_20__20_), .B(raddr2_0_bF_buf76_), .Y(_4960_) );
OAI21X1 OAI21X1_1916 ( .gnd(gnd), .vdd(vdd), .A(_1448_), .B(raddr2_0_bF_buf75_), .C(_4960_), .Y(_4961_) );
MUX2X1 MUX2X1_481 ( .gnd(gnd), .vdd(vdd), .A(_4961_), .B(_4959_), .S(raddr2_1_bF_buf11_), .Y(_4962_) );
NAND2X1 NAND2X1_948 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf3), .B(_4962_), .Y(_4963_) );
NAND2X1 NAND2X1_949 ( .gnd(gnd), .vdd(vdd), .A(regs_18__20_), .B(raddr2_0_bF_buf74_), .Y(_4964_) );
OAI21X1 OAI21X1_1917 ( .gnd(gnd), .vdd(vdd), .A(_1547_), .B(raddr2_0_bF_buf73_), .C(_4964_), .Y(_4965_) );
NAND2X1 NAND2X1_950 ( .gnd(gnd), .vdd(vdd), .A(regs_16__20_), .B(raddr2_0_bF_buf72_), .Y(_4966_) );
OAI21X1 OAI21X1_1918 ( .gnd(gnd), .vdd(vdd), .A(_1645_), .B(raddr2_0_bF_buf71_), .C(_4966_), .Y(_4967_) );
MUX2X1 MUX2X1_482 ( .gnd(gnd), .vdd(vdd), .A(_4967_), .B(_4965_), .S(raddr2_1_bF_buf10_), .Y(_4968_) );
AOI21X1 AOI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(raddr2_2_bF_buf4_), .B(_4968_), .C(_4033__bF_buf6), .Y(_4969_) );
OAI21X1 OAI21X1_1919 ( .gnd(gnd), .vdd(vdd), .A(_1183_), .B(raddr2_0_bF_buf70_), .C(raddr2_2_bF_buf3_), .Y(_4970_) );
AOI21X1 AOI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(regs_26__20_), .B(raddr2_0_bF_buf69_), .C(_4970_), .Y(_4971_) );
OAI21X1 OAI21X1_1920 ( .gnd(gnd), .vdd(vdd), .A(regs_30__20_), .B(raddr2_2_bF_buf2_), .C(_4038__bF_buf4), .Y(_4972_) );
OAI21X1 OAI21X1_1921 ( .gnd(gnd), .vdd(vdd), .A(_3468_), .B(raddr2_0_bF_buf68_), .C(raddr2_2_bF_buf1_), .Y(_4973_) );
AOI21X1 AOI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(regs_24__20_), .B(raddr2_0_bF_buf67_), .C(_4973_), .Y(_4974_) );
NOR2X1 NOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf66_), .B(_3462_), .Y(_4975_) );
NAND2X1 NAND2X1_951 ( .gnd(gnd), .vdd(vdd), .A(regs_28__20_), .B(raddr2_0_bF_buf65_), .Y(_4976_) );
NAND2X1 NAND2X1_952 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf2), .B(_4976_), .Y(_4977_) );
OAI21X1 OAI21X1_1922 ( .gnd(gnd), .vdd(vdd), .A(_4977_), .B(_4975_), .C(raddr2_1_bF_buf9_), .Y(_4978_) );
OAI22X1 OAI22X1_87 ( .gnd(gnd), .vdd(vdd), .A(_4971_), .B(_4972_), .C(_4978_), .D(_4974_), .Y(_4979_) );
AOI22X1 AOI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_4979_), .B(_4033__bF_buf5), .C(_4963_), .D(_4969_), .Y(_4980_) );
NAND2X1 NAND2X1_953 ( .gnd(gnd), .vdd(vdd), .A(regs_6__20_), .B(raddr2_0_bF_buf64_), .Y(_4981_) );
OAI21X1 OAI21X1_1923 ( .gnd(gnd), .vdd(vdd), .A(_2141_), .B(raddr2_0_bF_buf63_), .C(_4981_), .Y(_4982_) );
NAND2X1 NAND2X1_954 ( .gnd(gnd), .vdd(vdd), .A(regs_4__20_), .B(raddr2_0_bF_buf62_), .Y(_4983_) );
OAI21X1 OAI21X1_1924 ( .gnd(gnd), .vdd(vdd), .A(_3423_), .B(raddr2_0_bF_buf61_), .C(_4983_), .Y(_4984_) );
MUX2X1 MUX2X1_483 ( .gnd(gnd), .vdd(vdd), .A(_4984_), .B(_4982_), .S(raddr2_1_bF_buf8_), .Y(_4985_) );
NAND2X1 NAND2X1_955 ( .gnd(gnd), .vdd(vdd), .A(regs_2__20_), .B(raddr2_0_bF_buf60_), .Y(_4986_) );
OAI21X1 OAI21X1_1925 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .B(raddr2_0_bF_buf59_), .C(_4986_), .Y(_4987_) );
NAND2X1 NAND2X1_956 ( .gnd(gnd), .vdd(vdd), .A(regs_0__20_), .B(raddr2_0_bF_buf58_), .Y(_4988_) );
OAI21X1 OAI21X1_1926 ( .gnd(gnd), .vdd(vdd), .A(_3429_), .B(raddr2_0_bF_buf57_), .C(_4988_), .Y(_4989_) );
MUX2X1 MUX2X1_484 ( .gnd(gnd), .vdd(vdd), .A(_4989_), .B(_4987_), .S(raddr2_1_bF_buf7_), .Y(_4990_) );
MUX2X1 MUX2X1_485 ( .gnd(gnd), .vdd(vdd), .A(_4990_), .B(_4985_), .S(raddr2_2_bF_buf0_), .Y(_4991_) );
NAND2X1 NAND2X1_957 ( .gnd(gnd), .vdd(vdd), .A(regs_10__20_), .B(raddr2_0_bF_buf56_), .Y(_4992_) );
OAI21X1 OAI21X1_1927 ( .gnd(gnd), .vdd(vdd), .A(_1942_), .B(raddr2_0_bF_buf55_), .C(_4992_), .Y(_4993_) );
NAND2X1 NAND2X1_958 ( .gnd(gnd), .vdd(vdd), .A(regs_8__20_), .B(raddr2_0_bF_buf54_), .Y(_4994_) );
OAI21X1 OAI21X1_1928 ( .gnd(gnd), .vdd(vdd), .A(_2040_), .B(raddr2_0_bF_buf53_), .C(_4994_), .Y(_4995_) );
MUX2X1 MUX2X1_486 ( .gnd(gnd), .vdd(vdd), .A(_4995_), .B(_4993_), .S(raddr2_1_bF_buf6_), .Y(_4996_) );
NAND2X1 NAND2X1_959 ( .gnd(gnd), .vdd(vdd), .A(regs_14__20_), .B(raddr2_0_bF_buf52_), .Y(_4997_) );
OAI21X1 OAI21X1_1929 ( .gnd(gnd), .vdd(vdd), .A(_1745_), .B(raddr2_0_bF_buf51_), .C(_4997_), .Y(_4998_) );
NAND2X1 NAND2X1_960 ( .gnd(gnd), .vdd(vdd), .A(regs_12__20_), .B(raddr2_0_bF_buf50_), .Y(_4999_) );
OAI21X1 OAI21X1_1930 ( .gnd(gnd), .vdd(vdd), .A(_1843_), .B(raddr2_0_bF_buf49_), .C(_4999_), .Y(_5000_) );
MUX2X1 MUX2X1_487 ( .gnd(gnd), .vdd(vdd), .A(_5000_), .B(_4998_), .S(raddr2_1_bF_buf5_), .Y(_5001_) );
MUX2X1 MUX2X1_488 ( .gnd(gnd), .vdd(vdd), .A(_5001_), .B(_4996_), .S(_4036__bF_buf1), .Y(_5002_) );
MUX2X1 MUX2X1_489 ( .gnd(gnd), .vdd(vdd), .A(_5002_), .B(_4991_), .S(_4033__bF_buf4), .Y(_5003_) );
MUX2X1 MUX2X1_490 ( .gnd(gnd), .vdd(vdd), .A(_5003_), .B(_4980_), .S(raddr2_4_bF_buf4_), .Y(_5512__20_) );
OAI21X1 OAI21X1_1931 ( .gnd(gnd), .vdd(vdd), .A(_1450_), .B(raddr2_0_bF_buf48_), .C(raddr2_1_bF_buf4_), .Y(_5004_) );
AOI21X1 AOI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(regs_20__21_), .B(raddr2_0_bF_buf47_), .C(_5004_), .Y(_5005_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(regs_22__21_), .B(raddr2_0_bF_buf46_), .Y(_5006_) );
OAI21X1 OAI21X1_1932 ( .gnd(gnd), .vdd(vdd), .A(_1352_), .B(raddr2_0_bF_buf45_), .C(_4038__bF_buf3), .Y(_5007_) );
OAI21X1 OAI21X1_1933 ( .gnd(gnd), .vdd(vdd), .A(_5007_), .B(_5006_), .C(_4036__bF_buf0), .Y(_5008_) );
OAI21X1 OAI21X1_1934 ( .gnd(gnd), .vdd(vdd), .A(_1647_), .B(raddr2_0_bF_buf44_), .C(raddr2_1_bF_buf3_), .Y(_5009_) );
AOI21X1 AOI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(regs_16__21_), .B(raddr2_0_bF_buf43_), .C(_5009_), .Y(_5010_) );
NOR2X1 NOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf42_), .B(_1549_), .Y(_5011_) );
NAND2X1 NAND2X1_961 ( .gnd(gnd), .vdd(vdd), .A(regs_18__21_), .B(raddr2_0_bF_buf41_), .Y(_5012_) );
NAND2X1 NAND2X1_962 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf2), .B(_5012_), .Y(_5013_) );
OAI21X1 OAI21X1_1935 ( .gnd(gnd), .vdd(vdd), .A(_5013_), .B(_5011_), .C(raddr2_2_bF_buf10_), .Y(_5014_) );
OAI22X1 OAI22X1_88 ( .gnd(gnd), .vdd(vdd), .A(_5010_), .B(_5014_), .C(_5008_), .D(_5005_), .Y(_5015_) );
NAND2X1 NAND2X1_963 ( .gnd(gnd), .vdd(vdd), .A(regs_28__21_), .B(raddr2_0_bF_buf40_), .Y(_5016_) );
OAI21X1 OAI21X1_1936 ( .gnd(gnd), .vdd(vdd), .A(_3513_), .B(raddr2_0_bF_buf39_), .C(_5016_), .Y(_5017_) );
MUX2X1 MUX2X1_491 ( .gnd(gnd), .vdd(vdd), .A(_5017_), .B(regs_30__21_), .S(raddr2_1_bF_buf2_), .Y(_5018_) );
NAND2X1 NAND2X1_964 ( .gnd(gnd), .vdd(vdd), .A(regs_26__21_), .B(raddr2_0_bF_buf38_), .Y(_5019_) );
OAI21X1 OAI21X1_1937 ( .gnd(gnd), .vdd(vdd), .A(_1185_), .B(raddr2_0_bF_buf37_), .C(_5019_), .Y(_5020_) );
NAND2X1 NAND2X1_965 ( .gnd(gnd), .vdd(vdd), .A(regs_24__21_), .B(raddr2_0_bF_buf36_), .Y(_5021_) );
OAI21X1 OAI21X1_1938 ( .gnd(gnd), .vdd(vdd), .A(_3519_), .B(raddr2_0_bF_buf35_), .C(_5021_), .Y(_5022_) );
MUX2X1 MUX2X1_492 ( .gnd(gnd), .vdd(vdd), .A(_5022_), .B(_5020_), .S(raddr2_1_bF_buf1_), .Y(_5023_) );
MUX2X1 MUX2X1_493 ( .gnd(gnd), .vdd(vdd), .A(_5023_), .B(_5018_), .S(raddr2_2_bF_buf9_), .Y(_5024_) );
MUX2X1 MUX2X1_494 ( .gnd(gnd), .vdd(vdd), .A(_5024_), .B(_5015_), .S(_4033__bF_buf3), .Y(_5025_) );
NAND2X1 NAND2X1_966 ( .gnd(gnd), .vdd(vdd), .A(regs_6__21_), .B(raddr2_0_bF_buf34_), .Y(_5026_) );
OAI21X1 OAI21X1_1939 ( .gnd(gnd), .vdd(vdd), .A(_2143_), .B(raddr2_0_bF_buf33_), .C(_5026_), .Y(_5027_) );
NAND2X1 NAND2X1_967 ( .gnd(gnd), .vdd(vdd), .A(regs_4__21_), .B(raddr2_0_bF_buf32_), .Y(_5028_) );
OAI21X1 OAI21X1_1940 ( .gnd(gnd), .vdd(vdd), .A(_3474_), .B(raddr2_0_bF_buf31_), .C(_5028_), .Y(_5029_) );
MUX2X1 MUX2X1_495 ( .gnd(gnd), .vdd(vdd), .A(_5029_), .B(_5027_), .S(raddr2_1_bF_buf0_), .Y(_5030_) );
NAND2X1 NAND2X1_968 ( .gnd(gnd), .vdd(vdd), .A(regs_2__21_), .B(raddr2_0_bF_buf30_), .Y(_5031_) );
OAI21X1 OAI21X1_1941 ( .gnd(gnd), .vdd(vdd), .A(_3483_), .B(raddr2_0_bF_buf29_), .C(_5031_), .Y(_5032_) );
NAND2X1 NAND2X1_969 ( .gnd(gnd), .vdd(vdd), .A(regs_0__21_), .B(raddr2_0_bF_buf28_), .Y(_5033_) );
OAI21X1 OAI21X1_1942 ( .gnd(gnd), .vdd(vdd), .A(_3480_), .B(raddr2_0_bF_buf27_), .C(_5033_), .Y(_5034_) );
MUX2X1 MUX2X1_496 ( .gnd(gnd), .vdd(vdd), .A(_5034_), .B(_5032_), .S(raddr2_1_bF_buf14_bF_buf0_), .Y(_5035_) );
MUX2X1 MUX2X1_497 ( .gnd(gnd), .vdd(vdd), .A(_5035_), .B(_5030_), .S(raddr2_2_bF_buf8_), .Y(_5036_) );
NAND2X1 NAND2X1_970 ( .gnd(gnd), .vdd(vdd), .A(regs_14__21_), .B(raddr2_0_bF_buf26_), .Y(_5037_) );
OAI21X1 OAI21X1_1943 ( .gnd(gnd), .vdd(vdd), .A(_1747_), .B(raddr2_0_bF_buf25_), .C(_5037_), .Y(_5038_) );
NAND2X1 NAND2X1_971 ( .gnd(gnd), .vdd(vdd), .A(regs_12__21_), .B(raddr2_0_bF_buf24_), .Y(_5039_) );
OAI21X1 OAI21X1_1944 ( .gnd(gnd), .vdd(vdd), .A(_1845_), .B(raddr2_0_bF_buf23_), .C(_5039_), .Y(_5040_) );
MUX2X1 MUX2X1_498 ( .gnd(gnd), .vdd(vdd), .A(_5040_), .B(_5038_), .S(raddr2_1_bF_buf13_bF_buf0_), .Y(_5041_) );
NAND2X1 NAND2X1_972 ( .gnd(gnd), .vdd(vdd), .A(regs_10__21_), .B(raddr2_0_bF_buf22_), .Y(_5042_) );
OAI21X1 OAI21X1_1945 ( .gnd(gnd), .vdd(vdd), .A(_1944_), .B(raddr2_0_bF_buf21_), .C(_5042_), .Y(_5043_) );
NAND2X1 NAND2X1_973 ( .gnd(gnd), .vdd(vdd), .A(regs_8__21_), .B(raddr2_0_bF_buf20_), .Y(_5044_) );
OAI21X1 OAI21X1_1946 ( .gnd(gnd), .vdd(vdd), .A(_2042_), .B(raddr2_0_bF_buf19_), .C(_5044_), .Y(_5045_) );
MUX2X1 MUX2X1_499 ( .gnd(gnd), .vdd(vdd), .A(_5045_), .B(_5043_), .S(raddr2_1_bF_buf12_bF_buf0_), .Y(_5046_) );
MUX2X1 MUX2X1_500 ( .gnd(gnd), .vdd(vdd), .A(_5046_), .B(_5041_), .S(raddr2_2_bF_buf7_), .Y(_5047_) );
MUX2X1 MUX2X1_501 ( .gnd(gnd), .vdd(vdd), .A(_5047_), .B(_5036_), .S(_4033__bF_buf2), .Y(_5048_) );
MUX2X1 MUX2X1_502 ( .gnd(gnd), .vdd(vdd), .A(_5048_), .B(_5025_), .S(raddr2_4_bF_buf3_), .Y(_5512__21_) );
NAND2X1 NAND2X1_974 ( .gnd(gnd), .vdd(vdd), .A(regs_22__22_), .B(raddr2_0_bF_buf18_), .Y(_5049_) );
OAI21X1 OAI21X1_1947 ( .gnd(gnd), .vdd(vdd), .A(_1354_), .B(raddr2_0_bF_buf17_), .C(_5049_), .Y(_5050_) );
NAND2X1 NAND2X1_975 ( .gnd(gnd), .vdd(vdd), .A(regs_20__22_), .B(raddr2_0_bF_buf16_), .Y(_5051_) );
OAI21X1 OAI21X1_1948 ( .gnd(gnd), .vdd(vdd), .A(_1452_), .B(raddr2_0_bF_buf15_), .C(_5051_), .Y(_5052_) );
MUX2X1 MUX2X1_503 ( .gnd(gnd), .vdd(vdd), .A(_5052_), .B(_5050_), .S(raddr2_1_bF_buf11_), .Y(_5053_) );
NAND2X1 NAND2X1_976 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf8), .B(_5053_), .Y(_5054_) );
NAND2X1 NAND2X1_977 ( .gnd(gnd), .vdd(vdd), .A(regs_18__22_), .B(raddr2_0_bF_buf14_), .Y(_5055_) );
OAI21X1 OAI21X1_1949 ( .gnd(gnd), .vdd(vdd), .A(_1551_), .B(raddr2_0_bF_buf13_), .C(_5055_), .Y(_5056_) );
NAND2X1 NAND2X1_978 ( .gnd(gnd), .vdd(vdd), .A(regs_16__22_), .B(raddr2_0_bF_buf12_), .Y(_5057_) );
OAI21X1 OAI21X1_1950 ( .gnd(gnd), .vdd(vdd), .A(_1649_), .B(raddr2_0_bF_buf11_), .C(_5057_), .Y(_5058_) );
MUX2X1 MUX2X1_504 ( .gnd(gnd), .vdd(vdd), .A(_5058_), .B(_5056_), .S(raddr2_1_bF_buf10_), .Y(_5059_) );
AOI21X1 AOI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(raddr2_2_bF_buf6_), .B(_5059_), .C(_4033__bF_buf1), .Y(_5060_) );
OAI21X1 OAI21X1_1951 ( .gnd(gnd), .vdd(vdd), .A(_1187_), .B(raddr2_0_bF_buf10_), .C(raddr2_2_bF_buf5_), .Y(_5061_) );
AOI21X1 AOI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(regs_26__22_), .B(raddr2_0_bF_buf9_), .C(_5061_), .Y(_5062_) );
OAI21X1 OAI21X1_1952 ( .gnd(gnd), .vdd(vdd), .A(regs_30__22_), .B(raddr2_2_bF_buf4_), .C(_4038__bF_buf1), .Y(_5063_) );
OAI21X1 OAI21X1_1953 ( .gnd(gnd), .vdd(vdd), .A(_3543_), .B(raddr2_0_bF_buf8_), .C(raddr2_2_bF_buf3_), .Y(_5064_) );
AOI21X1 AOI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(regs_24__22_), .B(raddr2_0_bF_buf7_), .C(_5064_), .Y(_5065_) );
NOR2X1 NOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf6_), .B(_3537_), .Y(_5066_) );
NAND2X1 NAND2X1_979 ( .gnd(gnd), .vdd(vdd), .A(regs_28__22_), .B(raddr2_0_bF_buf5_), .Y(_5067_) );
NAND2X1 NAND2X1_980 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf7), .B(_5067_), .Y(_5068_) );
OAI21X1 OAI21X1_1954 ( .gnd(gnd), .vdd(vdd), .A(_5068_), .B(_5066_), .C(raddr2_1_bF_buf9_), .Y(_5069_) );
OAI22X1 OAI22X1_89 ( .gnd(gnd), .vdd(vdd), .A(_5062_), .B(_5063_), .C(_5069_), .D(_5065_), .Y(_5070_) );
AOI22X1 AOI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_5070_), .B(_4033__bF_buf0), .C(_5054_), .D(_5060_), .Y(_5071_) );
OAI21X1 OAI21X1_1955 ( .gnd(gnd), .vdd(vdd), .A(_3551_), .B(raddr2_0_bF_buf4_), .C(raddr2_1_bF_buf8_), .Y(_5072_) );
AOI21X1 AOI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(regs_4__22_), .B(raddr2_0_bF_buf3_), .C(_5072_), .Y(_5073_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(regs_6__22_), .B(raddr2_0_bF_buf2_), .Y(_5074_) );
OAI21X1 OAI21X1_1956 ( .gnd(gnd), .vdd(vdd), .A(_2145_), .B(raddr2_0_bF_buf1_), .C(_4038__bF_buf0), .Y(_5075_) );
OAI21X1 OAI21X1_1957 ( .gnd(gnd), .vdd(vdd), .A(_5075_), .B(_5074_), .C(_4036__bF_buf6), .Y(_5076_) );
OAI21X1 OAI21X1_1958 ( .gnd(gnd), .vdd(vdd), .A(_3558_), .B(raddr2_0_bF_buf0_), .C(raddr2_1_bF_buf7_), .Y(_5077_) );
AOI21X1 AOI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(regs_0__22_), .B(raddr2_0_bF_buf96_), .C(_5077_), .Y(_5078_) );
NOR2X1 NOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf95_), .B(_3555_), .Y(_5079_) );
NAND2X1 NAND2X1_981 ( .gnd(gnd), .vdd(vdd), .A(regs_2__22_), .B(raddr2_0_bF_buf94_), .Y(_5080_) );
NAND2X1 NAND2X1_982 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf8), .B(_5080_), .Y(_5081_) );
OAI21X1 OAI21X1_1959 ( .gnd(gnd), .vdd(vdd), .A(_5081_), .B(_5079_), .C(raddr2_2_bF_buf2_), .Y(_5082_) );
OAI22X1 OAI22X1_90 ( .gnd(gnd), .vdd(vdd), .A(_5078_), .B(_5082_), .C(_5076_), .D(_5073_), .Y(_5083_) );
NAND2X1 NAND2X1_983 ( .gnd(gnd), .vdd(vdd), .A(regs_10__22_), .B(raddr2_0_bF_buf93_), .Y(_5084_) );
OAI21X1 OAI21X1_1960 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(raddr2_0_bF_buf92_), .C(_5084_), .Y(_5085_) );
NAND2X1 NAND2X1_984 ( .gnd(gnd), .vdd(vdd), .A(regs_8__22_), .B(raddr2_0_bF_buf91_), .Y(_5086_) );
OAI21X1 OAI21X1_1961 ( .gnd(gnd), .vdd(vdd), .A(_2044_), .B(raddr2_0_bF_buf90_), .C(_5086_), .Y(_5087_) );
MUX2X1 MUX2X1_505 ( .gnd(gnd), .vdd(vdd), .A(_5087_), .B(_5085_), .S(raddr2_1_bF_buf6_), .Y(_5088_) );
NAND2X1 NAND2X1_985 ( .gnd(gnd), .vdd(vdd), .A(regs_14__22_), .B(raddr2_0_bF_buf89_), .Y(_5089_) );
OAI21X1 OAI21X1_1962 ( .gnd(gnd), .vdd(vdd), .A(_1749_), .B(raddr2_0_bF_buf88_), .C(_5089_), .Y(_5090_) );
NAND2X1 NAND2X1_986 ( .gnd(gnd), .vdd(vdd), .A(regs_12__22_), .B(raddr2_0_bF_buf87_), .Y(_5091_) );
OAI21X1 OAI21X1_1963 ( .gnd(gnd), .vdd(vdd), .A(_1847_), .B(raddr2_0_bF_buf86_), .C(_5091_), .Y(_5092_) );
MUX2X1 MUX2X1_506 ( .gnd(gnd), .vdd(vdd), .A(_5092_), .B(_5090_), .S(raddr2_1_bF_buf5_), .Y(_5093_) );
MUX2X1 MUX2X1_507 ( .gnd(gnd), .vdd(vdd), .A(_5093_), .B(_5088_), .S(_4036__bF_buf5), .Y(_5094_) );
MUX2X1 MUX2X1_508 ( .gnd(gnd), .vdd(vdd), .A(_5094_), .B(_5083_), .S(_4033__bF_buf7), .Y(_5095_) );
MUX2X1 MUX2X1_509 ( .gnd(gnd), .vdd(vdd), .A(_5095_), .B(_5071_), .S(raddr2_4_bF_buf2_), .Y(_5512__22_) );
OAI21X1 OAI21X1_1964 ( .gnd(gnd), .vdd(vdd), .A(_1454_), .B(raddr2_0_bF_buf85_), .C(raddr2_1_bF_buf4_), .Y(_5096_) );
AOI21X1 AOI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(regs_20__23_), .B(raddr2_0_bF_buf84_), .C(_5096_), .Y(_5097_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(regs_22__23_), .B(raddr2_0_bF_buf83_), .Y(_5098_) );
OAI21X1 OAI21X1_1965 ( .gnd(gnd), .vdd(vdd), .A(_1356_), .B(raddr2_0_bF_buf82_), .C(_4038__bF_buf7), .Y(_5099_) );
OAI21X1 OAI21X1_1966 ( .gnd(gnd), .vdd(vdd), .A(_5099_), .B(_5098_), .C(_4036__bF_buf4), .Y(_5100_) );
OAI21X1 OAI21X1_1967 ( .gnd(gnd), .vdd(vdd), .A(_1651_), .B(raddr2_0_bF_buf81_), .C(raddr2_1_bF_buf3_), .Y(_5101_) );
AOI21X1 AOI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(regs_16__23_), .B(raddr2_0_bF_buf80_), .C(_5101_), .Y(_5102_) );
NOR2X1 NOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf79_), .B(_1553_), .Y(_5103_) );
NAND2X1 NAND2X1_987 ( .gnd(gnd), .vdd(vdd), .A(regs_18__23_), .B(raddr2_0_bF_buf78_), .Y(_5104_) );
NAND2X1 NAND2X1_988 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf6), .B(_5104_), .Y(_5105_) );
OAI21X1 OAI21X1_1968 ( .gnd(gnd), .vdd(vdd), .A(_5105_), .B(_5103_), .C(raddr2_2_bF_buf1_), .Y(_5106_) );
OAI22X1 OAI22X1_91 ( .gnd(gnd), .vdd(vdd), .A(_5102_), .B(_5106_), .C(_5100_), .D(_5097_), .Y(_5107_) );
NAND2X1 NAND2X1_989 ( .gnd(gnd), .vdd(vdd), .A(regs_28__23_), .B(raddr2_0_bF_buf77_), .Y(_5108_) );
OAI21X1 OAI21X1_1969 ( .gnd(gnd), .vdd(vdd), .A(_3587_), .B(raddr2_0_bF_buf76_), .C(_5108_), .Y(_5109_) );
MUX2X1 MUX2X1_510 ( .gnd(gnd), .vdd(vdd), .A(_5109_), .B(regs_30__23_), .S(raddr2_1_bF_buf2_), .Y(_5110_) );
NAND2X1 NAND2X1_990 ( .gnd(gnd), .vdd(vdd), .A(regs_26__23_), .B(raddr2_0_bF_buf75_), .Y(_5111_) );
OAI21X1 OAI21X1_1970 ( .gnd(gnd), .vdd(vdd), .A(_1189_), .B(raddr2_0_bF_buf74_), .C(_5111_), .Y(_5112_) );
NAND2X1 NAND2X1_991 ( .gnd(gnd), .vdd(vdd), .A(regs_24__23_), .B(raddr2_0_bF_buf73_), .Y(_5113_) );
OAI21X1 OAI21X1_1971 ( .gnd(gnd), .vdd(vdd), .A(_3593_), .B(raddr2_0_bF_buf72_), .C(_5113_), .Y(_5114_) );
MUX2X1 MUX2X1_511 ( .gnd(gnd), .vdd(vdd), .A(_5114_), .B(_5112_), .S(raddr2_1_bF_buf1_), .Y(_5115_) );
MUX2X1 MUX2X1_512 ( .gnd(gnd), .vdd(vdd), .A(_5115_), .B(_5110_), .S(raddr2_2_bF_buf0_), .Y(_5116_) );
MUX2X1 MUX2X1_513 ( .gnd(gnd), .vdd(vdd), .A(_5116_), .B(_5107_), .S(_4033__bF_buf6), .Y(_5117_) );
NAND2X1 NAND2X1_992 ( .gnd(gnd), .vdd(vdd), .A(regs_6__23_), .B(raddr2_0_bF_buf71_), .Y(_5118_) );
OAI21X1 OAI21X1_1972 ( .gnd(gnd), .vdd(vdd), .A(_2147_), .B(raddr2_0_bF_buf70_), .C(_5118_), .Y(_5119_) );
NAND2X1 NAND2X1_993 ( .gnd(gnd), .vdd(vdd), .A(regs_4__23_), .B(raddr2_0_bF_buf69_), .Y(_5120_) );
OAI21X1 OAI21X1_1973 ( .gnd(gnd), .vdd(vdd), .A(_3601_), .B(raddr2_0_bF_buf68_), .C(_5120_), .Y(_5121_) );
MUX2X1 MUX2X1_514 ( .gnd(gnd), .vdd(vdd), .A(_5121_), .B(_5119_), .S(raddr2_1_bF_buf0_), .Y(_5122_) );
NAND2X1 NAND2X1_994 ( .gnd(gnd), .vdd(vdd), .A(regs_2__23_), .B(raddr2_0_bF_buf67_), .Y(_5123_) );
OAI21X1 OAI21X1_1974 ( .gnd(gnd), .vdd(vdd), .A(_3605_), .B(raddr2_0_bF_buf66_), .C(_5123_), .Y(_5124_) );
NAND2X1 NAND2X1_995 ( .gnd(gnd), .vdd(vdd), .A(regs_0__23_), .B(raddr2_0_bF_buf65_), .Y(_5125_) );
OAI21X1 OAI21X1_1975 ( .gnd(gnd), .vdd(vdd), .A(_3608_), .B(raddr2_0_bF_buf64_), .C(_5125_), .Y(_5126_) );
MUX2X1 MUX2X1_515 ( .gnd(gnd), .vdd(vdd), .A(_5126_), .B(_5124_), .S(raddr2_1_bF_buf14_bF_buf3_), .Y(_5127_) );
MUX2X1 MUX2X1_516 ( .gnd(gnd), .vdd(vdd), .A(_5127_), .B(_5122_), .S(raddr2_2_bF_buf10_), .Y(_5128_) );
NAND2X1 NAND2X1_996 ( .gnd(gnd), .vdd(vdd), .A(regs_10__23_), .B(raddr2_0_bF_buf63_), .Y(_5129_) );
OAI21X1 OAI21X1_1976 ( .gnd(gnd), .vdd(vdd), .A(_1948_), .B(raddr2_0_bF_buf62_), .C(_5129_), .Y(_5130_) );
NAND2X1 NAND2X1_997 ( .gnd(gnd), .vdd(vdd), .A(regs_8__23_), .B(raddr2_0_bF_buf61_), .Y(_5131_) );
OAI21X1 OAI21X1_1977 ( .gnd(gnd), .vdd(vdd), .A(_2046_), .B(raddr2_0_bF_buf60_), .C(_5131_), .Y(_5132_) );
MUX2X1 MUX2X1_517 ( .gnd(gnd), .vdd(vdd), .A(_5132_), .B(_5130_), .S(raddr2_1_bF_buf13_bF_buf3_), .Y(_5133_) );
NAND2X1 NAND2X1_998 ( .gnd(gnd), .vdd(vdd), .A(regs_14__23_), .B(raddr2_0_bF_buf59_), .Y(_5134_) );
OAI21X1 OAI21X1_1978 ( .gnd(gnd), .vdd(vdd), .A(_1751_), .B(raddr2_0_bF_buf58_), .C(_5134_), .Y(_5135_) );
NAND2X1 NAND2X1_999 ( .gnd(gnd), .vdd(vdd), .A(regs_12__23_), .B(raddr2_0_bF_buf57_), .Y(_5136_) );
OAI21X1 OAI21X1_1979 ( .gnd(gnd), .vdd(vdd), .A(_1849_), .B(raddr2_0_bF_buf56_), .C(_5136_), .Y(_5137_) );
MUX2X1 MUX2X1_518 ( .gnd(gnd), .vdd(vdd), .A(_5137_), .B(_5135_), .S(raddr2_1_bF_buf12_bF_buf3_), .Y(_5138_) );
MUX2X1 MUX2X1_519 ( .gnd(gnd), .vdd(vdd), .A(_5138_), .B(_5133_), .S(_4036__bF_buf3), .Y(_5139_) );
MUX2X1 MUX2X1_520 ( .gnd(gnd), .vdd(vdd), .A(_5139_), .B(_5128_), .S(_4033__bF_buf5), .Y(_5140_) );
MUX2X1 MUX2X1_521 ( .gnd(gnd), .vdd(vdd), .A(_5140_), .B(_5117_), .S(raddr2_4_bF_buf1_), .Y(_5512__23_) );
NAND2X1 NAND2X1_1000 ( .gnd(gnd), .vdd(vdd), .A(regs_22__24_), .B(raddr2_0_bF_buf55_), .Y(_5141_) );
OAI21X1 OAI21X1_1980 ( .gnd(gnd), .vdd(vdd), .A(_1358_), .B(raddr2_0_bF_buf54_), .C(_5141_), .Y(_5142_) );
NAND2X1 NAND2X1_1001 ( .gnd(gnd), .vdd(vdd), .A(regs_20__24_), .B(raddr2_0_bF_buf53_), .Y(_5143_) );
OAI21X1 OAI21X1_1981 ( .gnd(gnd), .vdd(vdd), .A(_1456_), .B(raddr2_0_bF_buf52_), .C(_5143_), .Y(_5144_) );
MUX2X1 MUX2X1_522 ( .gnd(gnd), .vdd(vdd), .A(_5144_), .B(_5142_), .S(raddr2_1_bF_buf11_), .Y(_5145_) );
NAND2X1 NAND2X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf2), .B(_5145_), .Y(_5146_) );
NAND2X1 NAND2X1_1003 ( .gnd(gnd), .vdd(vdd), .A(regs_18__24_), .B(raddr2_0_bF_buf51_), .Y(_5147_) );
OAI21X1 OAI21X1_1982 ( .gnd(gnd), .vdd(vdd), .A(_1555_), .B(raddr2_0_bF_buf50_), .C(_5147_), .Y(_5148_) );
NAND2X1 NAND2X1_1004 ( .gnd(gnd), .vdd(vdd), .A(regs_16__24_), .B(raddr2_0_bF_buf49_), .Y(_5149_) );
OAI21X1 OAI21X1_1983 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .B(raddr2_0_bF_buf48_), .C(_5149_), .Y(_5150_) );
MUX2X1 MUX2X1_523 ( .gnd(gnd), .vdd(vdd), .A(_5150_), .B(_5148_), .S(raddr2_1_bF_buf10_), .Y(_5151_) );
AOI21X1 AOI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(raddr2_2_bF_buf9_), .B(_5151_), .C(_4033__bF_buf4), .Y(_5152_) );
OAI21X1 OAI21X1_1984 ( .gnd(gnd), .vdd(vdd), .A(_1191_), .B(raddr2_0_bF_buf47_), .C(raddr2_2_bF_buf8_), .Y(_5153_) );
AOI21X1 AOI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(regs_26__24_), .B(raddr2_0_bF_buf46_), .C(_5153_), .Y(_5154_) );
OAI21X1 OAI21X1_1985 ( .gnd(gnd), .vdd(vdd), .A(regs_30__24_), .B(raddr2_2_bF_buf7_), .C(_4038__bF_buf5), .Y(_5155_) );
OAI21X1 OAI21X1_1986 ( .gnd(gnd), .vdd(vdd), .A(_3643_), .B(raddr2_0_bF_buf45_), .C(raddr2_2_bF_buf6_), .Y(_5156_) );
AOI21X1 AOI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(regs_24__24_), .B(raddr2_0_bF_buf44_), .C(_5156_), .Y(_5157_) );
NOR2X1 NOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf43_), .B(_3637_), .Y(_5158_) );
NAND2X1 NAND2X1_1005 ( .gnd(gnd), .vdd(vdd), .A(regs_28__24_), .B(raddr2_0_bF_buf42_), .Y(_5159_) );
NAND2X1 NAND2X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf1), .B(_5159_), .Y(_5160_) );
OAI21X1 OAI21X1_1987 ( .gnd(gnd), .vdd(vdd), .A(_5160_), .B(_5158_), .C(raddr2_1_bF_buf9_), .Y(_5161_) );
OAI22X1 OAI22X1_92 ( .gnd(gnd), .vdd(vdd), .A(_5154_), .B(_5155_), .C(_5161_), .D(_5157_), .Y(_5162_) );
AOI22X1 AOI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_5162_), .B(_4033__bF_buf3), .C(_5146_), .D(_5152_), .Y(_5163_) );
OAI21X1 OAI21X1_1988 ( .gnd(gnd), .vdd(vdd), .A(_3651_), .B(raddr2_0_bF_buf41_), .C(raddr2_1_bF_buf8_), .Y(_5164_) );
AOI21X1 AOI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(regs_4__24_), .B(raddr2_0_bF_buf40_), .C(_5164_), .Y(_5165_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(regs_6__24_), .B(raddr2_0_bF_buf39_), .Y(_5166_) );
OAI21X1 OAI21X1_1989 ( .gnd(gnd), .vdd(vdd), .A(_2149_), .B(raddr2_0_bF_buf38_), .C(_4038__bF_buf4), .Y(_5167_) );
OAI21X1 OAI21X1_1990 ( .gnd(gnd), .vdd(vdd), .A(_5167_), .B(_5166_), .C(_4036__bF_buf0), .Y(_5168_) );
OAI21X1 OAI21X1_1991 ( .gnd(gnd), .vdd(vdd), .A(_3658_), .B(raddr2_0_bF_buf37_), .C(raddr2_1_bF_buf7_), .Y(_5169_) );
AOI21X1 AOI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(regs_0__24_), .B(raddr2_0_bF_buf36_), .C(_5169_), .Y(_5170_) );
NOR2X1 NOR2X1_234 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf35_), .B(_3655_), .Y(_5171_) );
NAND2X1 NAND2X1_1007 ( .gnd(gnd), .vdd(vdd), .A(regs_2__24_), .B(raddr2_0_bF_buf34_), .Y(_5172_) );
NAND2X1 NAND2X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf3), .B(_5172_), .Y(_5173_) );
OAI21X1 OAI21X1_1992 ( .gnd(gnd), .vdd(vdd), .A(_5173_), .B(_5171_), .C(raddr2_2_bF_buf5_), .Y(_5174_) );
OAI22X1 OAI22X1_93 ( .gnd(gnd), .vdd(vdd), .A(_5170_), .B(_5174_), .C(_5168_), .D(_5165_), .Y(_5175_) );
NAND2X1 NAND2X1_1009 ( .gnd(gnd), .vdd(vdd), .A(regs_10__24_), .B(raddr2_0_bF_buf33_), .Y(_5176_) );
OAI21X1 OAI21X1_1993 ( .gnd(gnd), .vdd(vdd), .A(_1950_), .B(raddr2_0_bF_buf32_), .C(_5176_), .Y(_5177_) );
NAND2X1 NAND2X1_1010 ( .gnd(gnd), .vdd(vdd), .A(regs_8__24_), .B(raddr2_0_bF_buf31_), .Y(_5178_) );
OAI21X1 OAI21X1_1994 ( .gnd(gnd), .vdd(vdd), .A(_2048_), .B(raddr2_0_bF_buf30_), .C(_5178_), .Y(_5179_) );
MUX2X1 MUX2X1_524 ( .gnd(gnd), .vdd(vdd), .A(_5179_), .B(_5177_), .S(raddr2_1_bF_buf6_), .Y(_5180_) );
NAND2X1 NAND2X1_1011 ( .gnd(gnd), .vdd(vdd), .A(regs_14__24_), .B(raddr2_0_bF_buf29_), .Y(_5181_) );
OAI21X1 OAI21X1_1995 ( .gnd(gnd), .vdd(vdd), .A(_1753_), .B(raddr2_0_bF_buf28_), .C(_5181_), .Y(_5182_) );
NAND2X1 NAND2X1_1012 ( .gnd(gnd), .vdd(vdd), .A(regs_12__24_), .B(raddr2_0_bF_buf27_), .Y(_5183_) );
OAI21X1 OAI21X1_1996 ( .gnd(gnd), .vdd(vdd), .A(_1851_), .B(raddr2_0_bF_buf26_), .C(_5183_), .Y(_5184_) );
MUX2X1 MUX2X1_525 ( .gnd(gnd), .vdd(vdd), .A(_5184_), .B(_5182_), .S(raddr2_1_bF_buf5_), .Y(_5185_) );
MUX2X1 MUX2X1_526 ( .gnd(gnd), .vdd(vdd), .A(_5185_), .B(_5180_), .S(_4036__bF_buf8), .Y(_5186_) );
MUX2X1 MUX2X1_527 ( .gnd(gnd), .vdd(vdd), .A(_5186_), .B(_5175_), .S(_4033__bF_buf2), .Y(_5187_) );
MUX2X1 MUX2X1_528 ( .gnd(gnd), .vdd(vdd), .A(_5187_), .B(_5163_), .S(raddr2_4_bF_buf0_), .Y(_5512__24_) );
NAND2X1 NAND2X1_1013 ( .gnd(gnd), .vdd(vdd), .A(regs_22__25_), .B(raddr2_0_bF_buf25_), .Y(_5188_) );
OAI21X1 OAI21X1_1997 ( .gnd(gnd), .vdd(vdd), .A(_1360_), .B(raddr2_0_bF_buf24_), .C(_5188_), .Y(_5189_) );
NAND2X1 NAND2X1_1014 ( .gnd(gnd), .vdd(vdd), .A(regs_20__25_), .B(raddr2_0_bF_buf23_), .Y(_5190_) );
OAI21X1 OAI21X1_1998 ( .gnd(gnd), .vdd(vdd), .A(_1458_), .B(raddr2_0_bF_buf22_), .C(_5190_), .Y(_5191_) );
MUX2X1 MUX2X1_529 ( .gnd(gnd), .vdd(vdd), .A(_5191_), .B(_5189_), .S(raddr2_1_bF_buf4_), .Y(_5192_) );
NAND2X1 NAND2X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf7), .B(_5192_), .Y(_5193_) );
NAND2X1 NAND2X1_1016 ( .gnd(gnd), .vdd(vdd), .A(regs_18__25_), .B(raddr2_0_bF_buf21_), .Y(_5194_) );
OAI21X1 OAI21X1_1999 ( .gnd(gnd), .vdd(vdd), .A(_1557_), .B(raddr2_0_bF_buf20_), .C(_5194_), .Y(_5195_) );
NAND2X1 NAND2X1_1017 ( .gnd(gnd), .vdd(vdd), .A(regs_16__25_), .B(raddr2_0_bF_buf19_), .Y(_5196_) );
OAI21X1 OAI21X1_2000 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .B(raddr2_0_bF_buf18_), .C(_5196_), .Y(_5197_) );
MUX2X1 MUX2X1_530 ( .gnd(gnd), .vdd(vdd), .A(_5197_), .B(_5195_), .S(raddr2_1_bF_buf3_), .Y(_5198_) );
AOI21X1 AOI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(raddr2_2_bF_buf4_), .B(_5198_), .C(_4033__bF_buf1), .Y(_5199_) );
OAI21X1 OAI21X1_2001 ( .gnd(gnd), .vdd(vdd), .A(_1193_), .B(raddr2_0_bF_buf17_), .C(raddr2_2_bF_buf3_), .Y(_5200_) );
AOI21X1 AOI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(regs_26__25_), .B(raddr2_0_bF_buf16_), .C(_5200_), .Y(_5201_) );
OAI21X1 OAI21X1_2002 ( .gnd(gnd), .vdd(vdd), .A(regs_30__25_), .B(raddr2_2_bF_buf2_), .C(_4038__bF_buf2), .Y(_5202_) );
OAI21X1 OAI21X1_2003 ( .gnd(gnd), .vdd(vdd), .A(_3720_), .B(raddr2_0_bF_buf15_), .C(raddr2_2_bF_buf1_), .Y(_5203_) );
AOI21X1 AOI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(regs_24__25_), .B(raddr2_0_bF_buf14_), .C(_5203_), .Y(_5204_) );
NOR2X1 NOR2X1_235 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf13_), .B(_3714_), .Y(_5205_) );
NAND2X1 NAND2X1_1018 ( .gnd(gnd), .vdd(vdd), .A(regs_28__25_), .B(raddr2_0_bF_buf12_), .Y(_5206_) );
NAND2X1 NAND2X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf6), .B(_5206_), .Y(_5207_) );
OAI21X1 OAI21X1_2004 ( .gnd(gnd), .vdd(vdd), .A(_5207_), .B(_5205_), .C(raddr2_1_bF_buf2_), .Y(_5208_) );
OAI22X1 OAI22X1_94 ( .gnd(gnd), .vdd(vdd), .A(_5201_), .B(_5202_), .C(_5208_), .D(_5204_), .Y(_5209_) );
AOI22X1 AOI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_5209_), .B(_4033__bF_buf0), .C(_5193_), .D(_5199_), .Y(_5210_) );
NAND2X1 NAND2X1_1020 ( .gnd(gnd), .vdd(vdd), .A(regs_6__25_), .B(raddr2_0_bF_buf11_), .Y(_5211_) );
OAI21X1 OAI21X1_2005 ( .gnd(gnd), .vdd(vdd), .A(_2151_), .B(raddr2_0_bF_buf10_), .C(_5211_), .Y(_5212_) );
NAND2X1 NAND2X1_1021 ( .gnd(gnd), .vdd(vdd), .A(regs_4__25_), .B(raddr2_0_bF_buf9_), .Y(_5213_) );
OAI21X1 OAI21X1_2006 ( .gnd(gnd), .vdd(vdd), .A(_3675_), .B(raddr2_0_bF_buf8_), .C(_5213_), .Y(_5214_) );
MUX2X1 MUX2X1_531 ( .gnd(gnd), .vdd(vdd), .A(_5214_), .B(_5212_), .S(raddr2_1_bF_buf1_), .Y(_5215_) );
NAND2X1 NAND2X1_1022 ( .gnd(gnd), .vdd(vdd), .A(regs_2__25_), .B(raddr2_0_bF_buf7_), .Y(_5216_) );
OAI21X1 OAI21X1_2007 ( .gnd(gnd), .vdd(vdd), .A(_3684_), .B(raddr2_0_bF_buf6_), .C(_5216_), .Y(_5217_) );
NAND2X1 NAND2X1_1023 ( .gnd(gnd), .vdd(vdd), .A(regs_0__25_), .B(raddr2_0_bF_buf5_), .Y(_5218_) );
OAI21X1 OAI21X1_2008 ( .gnd(gnd), .vdd(vdd), .A(_3681_), .B(raddr2_0_bF_buf4_), .C(_5218_), .Y(_5219_) );
MUX2X1 MUX2X1_532 ( .gnd(gnd), .vdd(vdd), .A(_5219_), .B(_5217_), .S(raddr2_1_bF_buf0_), .Y(_5220_) );
MUX2X1 MUX2X1_533 ( .gnd(gnd), .vdd(vdd), .A(_5220_), .B(_5215_), .S(raddr2_2_bF_buf0_), .Y(_5221_) );
NAND2X1 NAND2X1_1024 ( .gnd(gnd), .vdd(vdd), .A(regs_14__25_), .B(raddr2_0_bF_buf3_), .Y(_5222_) );
OAI21X1 OAI21X1_2009 ( .gnd(gnd), .vdd(vdd), .A(_1755_), .B(raddr2_0_bF_buf2_), .C(_5222_), .Y(_5223_) );
NAND2X1 NAND2X1_1025 ( .gnd(gnd), .vdd(vdd), .A(regs_12__25_), .B(raddr2_0_bF_buf1_), .Y(_5224_) );
OAI21X1 OAI21X1_2010 ( .gnd(gnd), .vdd(vdd), .A(_1853_), .B(raddr2_0_bF_buf0_), .C(_5224_), .Y(_5225_) );
MUX2X1 MUX2X1_534 ( .gnd(gnd), .vdd(vdd), .A(_5225_), .B(_5223_), .S(raddr2_1_bF_buf14_bF_buf2_), .Y(_5226_) );
NAND2X1 NAND2X1_1026 ( .gnd(gnd), .vdd(vdd), .A(regs_10__25_), .B(raddr2_0_bF_buf96_), .Y(_5227_) );
OAI21X1 OAI21X1_2011 ( .gnd(gnd), .vdd(vdd), .A(_1952_), .B(raddr2_0_bF_buf95_), .C(_5227_), .Y(_5228_) );
NAND2X1 NAND2X1_1027 ( .gnd(gnd), .vdd(vdd), .A(regs_8__25_), .B(raddr2_0_bF_buf94_), .Y(_5229_) );
OAI21X1 OAI21X1_2012 ( .gnd(gnd), .vdd(vdd), .A(_2050_), .B(raddr2_0_bF_buf93_), .C(_5229_), .Y(_5230_) );
MUX2X1 MUX2X1_535 ( .gnd(gnd), .vdd(vdd), .A(_5230_), .B(_5228_), .S(raddr2_1_bF_buf13_bF_buf2_), .Y(_5231_) );
MUX2X1 MUX2X1_536 ( .gnd(gnd), .vdd(vdd), .A(_5231_), .B(_5226_), .S(raddr2_2_bF_buf10_), .Y(_5232_) );
MUX2X1 MUX2X1_537 ( .gnd(gnd), .vdd(vdd), .A(_5232_), .B(_5221_), .S(_4033__bF_buf7), .Y(_5233_) );
MUX2X1 MUX2X1_538 ( .gnd(gnd), .vdd(vdd), .A(_5233_), .B(_5210_), .S(raddr2_4_bF_buf4_), .Y(_5512__25_) );
OAI21X1 OAI21X1_2013 ( .gnd(gnd), .vdd(vdd), .A(_3726_), .B(raddr2_0_bF_buf92_), .C(raddr2_1_bF_buf12_bF_buf2_), .Y(_5234_) );
AOI21X1 AOI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(regs_4__26_), .B(raddr2_0_bF_buf91_), .C(_5234_), .Y(_5235_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(regs_6__26_), .B(raddr2_0_bF_buf90_), .Y(_5236_) );
OAI21X1 OAI21X1_2014 ( .gnd(gnd), .vdd(vdd), .A(_2153_), .B(raddr2_0_bF_buf89_), .C(_4038__bF_buf1), .Y(_5237_) );
OAI21X1 OAI21X1_2015 ( .gnd(gnd), .vdd(vdd), .A(_5237_), .B(_5236_), .C(_4036__bF_buf5), .Y(_5238_) );
OAI21X1 OAI21X1_2016 ( .gnd(gnd), .vdd(vdd), .A(_3732_), .B(raddr2_0_bF_buf88_), .C(raddr2_1_bF_buf11_), .Y(_5239_) );
AOI21X1 AOI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(regs_0__26_), .B(raddr2_0_bF_buf87_), .C(_5239_), .Y(_5240_) );
NOR2X1 NOR2X1_236 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf86_), .B(_3735_), .Y(_5241_) );
NAND2X1 NAND2X1_1028 ( .gnd(gnd), .vdd(vdd), .A(regs_2__26_), .B(raddr2_0_bF_buf85_), .Y(_5242_) );
NAND2X1 NAND2X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf0), .B(_5242_), .Y(_5243_) );
OAI21X1 OAI21X1_2017 ( .gnd(gnd), .vdd(vdd), .A(_5243_), .B(_5241_), .C(raddr2_2_bF_buf9_), .Y(_5244_) );
OAI22X1 OAI22X1_95 ( .gnd(gnd), .vdd(vdd), .A(_5240_), .B(_5244_), .C(_5238_), .D(_5235_), .Y(_5245_) );
NAND2X1 NAND2X1_1030 ( .gnd(gnd), .vdd(vdd), .A(regs_10__26_), .B(raddr2_0_bF_buf84_), .Y(_5246_) );
OAI21X1 OAI21X1_2018 ( .gnd(gnd), .vdd(vdd), .A(_1954_), .B(raddr2_0_bF_buf83_), .C(_5246_), .Y(_5247_) );
NAND2X1 NAND2X1_1031 ( .gnd(gnd), .vdd(vdd), .A(regs_8__26_), .B(raddr2_0_bF_buf82_), .Y(_5248_) );
OAI21X1 OAI21X1_2019 ( .gnd(gnd), .vdd(vdd), .A(_2052_), .B(raddr2_0_bF_buf81_), .C(_5248_), .Y(_5249_) );
MUX2X1 MUX2X1_539 ( .gnd(gnd), .vdd(vdd), .A(_5249_), .B(_5247_), .S(raddr2_1_bF_buf10_), .Y(_5250_) );
NAND2X1 NAND2X1_1032 ( .gnd(gnd), .vdd(vdd), .A(regs_14__26_), .B(raddr2_0_bF_buf80_), .Y(_5251_) );
OAI21X1 OAI21X1_2020 ( .gnd(gnd), .vdd(vdd), .A(_1757_), .B(raddr2_0_bF_buf79_), .C(_5251_), .Y(_5252_) );
NAND2X1 NAND2X1_1033 ( .gnd(gnd), .vdd(vdd), .A(regs_12__26_), .B(raddr2_0_bF_buf78_), .Y(_5253_) );
OAI21X1 OAI21X1_2021 ( .gnd(gnd), .vdd(vdd), .A(_1855_), .B(raddr2_0_bF_buf77_), .C(_5253_), .Y(_5254_) );
MUX2X1 MUX2X1_540 ( .gnd(gnd), .vdd(vdd), .A(_5254_), .B(_5252_), .S(raddr2_1_bF_buf9_), .Y(_5255_) );
MUX2X1 MUX2X1_541 ( .gnd(gnd), .vdd(vdd), .A(_5255_), .B(_5250_), .S(_4036__bF_buf4), .Y(_5256_) );
MUX2X1 MUX2X1_542 ( .gnd(gnd), .vdd(vdd), .A(_5256_), .B(_5245_), .S(_4033__bF_buf6), .Y(_5257_) );
OAI21X1 OAI21X1_2022 ( .gnd(gnd), .vdd(vdd), .A(_1657_), .B(raddr2_0_bF_buf76_), .C(raddr2_1_bF_buf8_), .Y(_5258_) );
AOI21X1 AOI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(regs_16__26_), .B(raddr2_0_bF_buf75_), .C(_5258_), .Y(_5259_) );
NOR2X1 NOR2X1_237 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf74_), .B(_1559_), .Y(_5260_) );
NAND2X1 NAND2X1_1034 ( .gnd(gnd), .vdd(vdd), .A(regs_18__26_), .B(raddr2_0_bF_buf73_), .Y(_5261_) );
NAND2X1 NAND2X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf8), .B(_5261_), .Y(_5262_) );
OAI21X1 OAI21X1_2023 ( .gnd(gnd), .vdd(vdd), .A(_5262_), .B(_5260_), .C(raddr2_2_bF_buf8_), .Y(_5263_) );
OAI21X1 OAI21X1_2024 ( .gnd(gnd), .vdd(vdd), .A(_1460_), .B(raddr2_0_bF_buf72_), .C(raddr2_1_bF_buf7_), .Y(_5264_) );
AOI21X1 AOI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(regs_20__26_), .B(raddr2_0_bF_buf71_), .C(_5264_), .Y(_5265_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(regs_22__26_), .B(raddr2_0_bF_buf70_), .Y(_5266_) );
OAI21X1 OAI21X1_2025 ( .gnd(gnd), .vdd(vdd), .A(_1362_), .B(raddr2_0_bF_buf69_), .C(_4038__bF_buf7), .Y(_5267_) );
OAI21X1 OAI21X1_2026 ( .gnd(gnd), .vdd(vdd), .A(_5267_), .B(_5266_), .C(_4036__bF_buf3), .Y(_5268_) );
OAI22X1 OAI22X1_96 ( .gnd(gnd), .vdd(vdd), .A(_5259_), .B(_5263_), .C(_5268_), .D(_5265_), .Y(_5269_) );
NAND2X1 NAND2X1_1036 ( .gnd(gnd), .vdd(vdd), .A(regs_28__26_), .B(raddr2_0_bF_buf68_), .Y(_5270_) );
OAI21X1 OAI21X1_2027 ( .gnd(gnd), .vdd(vdd), .A(_3765_), .B(raddr2_0_bF_buf67_), .C(_5270_), .Y(_5271_) );
MUX2X1 MUX2X1_543 ( .gnd(gnd), .vdd(vdd), .A(_5271_), .B(regs_30__26_), .S(raddr2_1_bF_buf6_), .Y(_5272_) );
NAND2X1 NAND2X1_1037 ( .gnd(gnd), .vdd(vdd), .A(regs_26__26_), .B(raddr2_0_bF_buf66_), .Y(_5273_) );
OAI21X1 OAI21X1_2028 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(raddr2_0_bF_buf65_), .C(_5273_), .Y(_5274_) );
NAND2X1 NAND2X1_1038 ( .gnd(gnd), .vdd(vdd), .A(regs_24__26_), .B(raddr2_0_bF_buf64_), .Y(_5275_) );
OAI21X1 OAI21X1_2029 ( .gnd(gnd), .vdd(vdd), .A(_3771_), .B(raddr2_0_bF_buf63_), .C(_5275_), .Y(_5276_) );
MUX2X1 MUX2X1_544 ( .gnd(gnd), .vdd(vdd), .A(_5276_), .B(_5274_), .S(raddr2_1_bF_buf5_), .Y(_5277_) );
MUX2X1 MUX2X1_545 ( .gnd(gnd), .vdd(vdd), .A(_5277_), .B(_5272_), .S(raddr2_2_bF_buf7_), .Y(_5278_) );
MUX2X1 MUX2X1_546 ( .gnd(gnd), .vdd(vdd), .A(_5278_), .B(_5269_), .S(_4033__bF_buf5), .Y(_5279_) );
MUX2X1 MUX2X1_547 ( .gnd(gnd), .vdd(vdd), .A(_5257_), .B(_5279_), .S(raddr2_4_bF_buf3_), .Y(_5512__26_) );
OAI21X1 OAI21X1_2030 ( .gnd(gnd), .vdd(vdd), .A(_1462_), .B(raddr2_0_bF_buf62_), .C(raddr2_1_bF_buf4_), .Y(_5280_) );
AOI21X1 AOI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(regs_20__27_), .B(raddr2_0_bF_buf61_), .C(_5280_), .Y(_5281_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(regs_22__27_), .B(raddr2_0_bF_buf60_), .Y(_5282_) );
OAI21X1 OAI21X1_2031 ( .gnd(gnd), .vdd(vdd), .A(_1364_), .B(raddr2_0_bF_buf59_), .C(_4038__bF_buf6), .Y(_5283_) );
OAI21X1 OAI21X1_2032 ( .gnd(gnd), .vdd(vdd), .A(_5283_), .B(_5282_), .C(_4036__bF_buf2), .Y(_5284_) );
OAI21X1 OAI21X1_2033 ( .gnd(gnd), .vdd(vdd), .A(_1659_), .B(raddr2_0_bF_buf58_), .C(raddr2_1_bF_buf3_), .Y(_5285_) );
AOI21X1 AOI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(regs_16__27_), .B(raddr2_0_bF_buf57_), .C(_5285_), .Y(_5286_) );
NOR2X1 NOR2X1_238 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf56_), .B(_1561_), .Y(_5287_) );
NAND2X1 NAND2X1_1039 ( .gnd(gnd), .vdd(vdd), .A(regs_18__27_), .B(raddr2_0_bF_buf55_), .Y(_5288_) );
NAND2X1 NAND2X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf5), .B(_5288_), .Y(_5289_) );
OAI21X1 OAI21X1_2034 ( .gnd(gnd), .vdd(vdd), .A(_5289_), .B(_5287_), .C(raddr2_2_bF_buf6_), .Y(_5290_) );
OAI22X1 OAI22X1_97 ( .gnd(gnd), .vdd(vdd), .A(_5286_), .B(_5290_), .C(_5284_), .D(_5281_), .Y(_5291_) );
NAND2X1 NAND2X1_1041 ( .gnd(gnd), .vdd(vdd), .A(regs_28__27_), .B(raddr2_0_bF_buf54_), .Y(_5292_) );
OAI21X1 OAI21X1_2035 ( .gnd(gnd), .vdd(vdd), .A(_3795_), .B(raddr2_0_bF_buf53_), .C(_5292_), .Y(_5293_) );
MUX2X1 MUX2X1_548 ( .gnd(gnd), .vdd(vdd), .A(_5293_), .B(regs_30__27_), .S(raddr2_1_bF_buf2_), .Y(_5294_) );
NAND2X1 NAND2X1_1042 ( .gnd(gnd), .vdd(vdd), .A(regs_26__27_), .B(raddr2_0_bF_buf52_), .Y(_5295_) );
OAI21X1 OAI21X1_2036 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(raddr2_0_bF_buf51_), .C(_5295_), .Y(_5296_) );
NAND2X1 NAND2X1_1043 ( .gnd(gnd), .vdd(vdd), .A(regs_24__27_), .B(raddr2_0_bF_buf50_), .Y(_5297_) );
OAI21X1 OAI21X1_2037 ( .gnd(gnd), .vdd(vdd), .A(_3792_), .B(raddr2_0_bF_buf49_), .C(_5297_), .Y(_5298_) );
MUX2X1 MUX2X1_549 ( .gnd(gnd), .vdd(vdd), .A(_5298_), .B(_5296_), .S(raddr2_1_bF_buf1_), .Y(_5299_) );
MUX2X1 MUX2X1_550 ( .gnd(gnd), .vdd(vdd), .A(_5299_), .B(_5294_), .S(raddr2_2_bF_buf5_), .Y(_5300_) );
MUX2X1 MUX2X1_551 ( .gnd(gnd), .vdd(vdd), .A(_5300_), .B(_5291_), .S(_4033__bF_buf4), .Y(_5301_) );
NAND2X1 NAND2X1_1044 ( .gnd(gnd), .vdd(vdd), .A(regs_6__27_), .B(raddr2_0_bF_buf48_), .Y(_5302_) );
OAI21X1 OAI21X1_2038 ( .gnd(gnd), .vdd(vdd), .A(_2155_), .B(raddr2_0_bF_buf47_), .C(_5302_), .Y(_5303_) );
NAND2X1 NAND2X1_1045 ( .gnd(gnd), .vdd(vdd), .A(regs_4__27_), .B(raddr2_0_bF_buf46_), .Y(_5304_) );
OAI21X1 OAI21X1_2039 ( .gnd(gnd), .vdd(vdd), .A(_3804_), .B(raddr2_0_bF_buf45_), .C(_5304_), .Y(_5305_) );
MUX2X1 MUX2X1_552 ( .gnd(gnd), .vdd(vdd), .A(_5305_), .B(_5303_), .S(raddr2_1_bF_buf0_), .Y(_5306_) );
NAND2X1 NAND2X1_1046 ( .gnd(gnd), .vdd(vdd), .A(regs_2__27_), .B(raddr2_0_bF_buf44_), .Y(_5307_) );
OAI21X1 OAI21X1_2040 ( .gnd(gnd), .vdd(vdd), .A(_3808_), .B(raddr2_0_bF_buf43_), .C(_5307_), .Y(_5308_) );
NAND2X1 NAND2X1_1047 ( .gnd(gnd), .vdd(vdd), .A(regs_0__27_), .B(raddr2_0_bF_buf42_), .Y(_5309_) );
OAI21X1 OAI21X1_2041 ( .gnd(gnd), .vdd(vdd), .A(_3811_), .B(raddr2_0_bF_buf41_), .C(_5309_), .Y(_5310_) );
MUX2X1 MUX2X1_553 ( .gnd(gnd), .vdd(vdd), .A(_5310_), .B(_5308_), .S(raddr2_1_bF_buf14_bF_buf1_), .Y(_5311_) );
MUX2X1 MUX2X1_554 ( .gnd(gnd), .vdd(vdd), .A(_5311_), .B(_5306_), .S(raddr2_2_bF_buf4_), .Y(_5312_) );
NAND2X1 NAND2X1_1048 ( .gnd(gnd), .vdd(vdd), .A(regs_10__27_), .B(raddr2_0_bF_buf40_), .Y(_5313_) );
OAI21X1 OAI21X1_2042 ( .gnd(gnd), .vdd(vdd), .A(_1956_), .B(raddr2_0_bF_buf39_), .C(_5313_), .Y(_5314_) );
NAND2X1 NAND2X1_1049 ( .gnd(gnd), .vdd(vdd), .A(regs_8__27_), .B(raddr2_0_bF_buf38_), .Y(_5315_) );
OAI21X1 OAI21X1_2043 ( .gnd(gnd), .vdd(vdd), .A(_2054_), .B(raddr2_0_bF_buf37_), .C(_5315_), .Y(_5316_) );
MUX2X1 MUX2X1_555 ( .gnd(gnd), .vdd(vdd), .A(_5316_), .B(_5314_), .S(raddr2_1_bF_buf13_bF_buf1_), .Y(_5317_) );
NAND2X1 NAND2X1_1050 ( .gnd(gnd), .vdd(vdd), .A(regs_14__27_), .B(raddr2_0_bF_buf36_), .Y(_5318_) );
OAI21X1 OAI21X1_2044 ( .gnd(gnd), .vdd(vdd), .A(_1759_), .B(raddr2_0_bF_buf35_), .C(_5318_), .Y(_5319_) );
NAND2X1 NAND2X1_1051 ( .gnd(gnd), .vdd(vdd), .A(regs_12__27_), .B(raddr2_0_bF_buf34_), .Y(_5320_) );
OAI21X1 OAI21X1_2045 ( .gnd(gnd), .vdd(vdd), .A(_1857_), .B(raddr2_0_bF_buf33_), .C(_5320_), .Y(_5321_) );
MUX2X1 MUX2X1_556 ( .gnd(gnd), .vdd(vdd), .A(_5321_), .B(_5319_), .S(raddr2_1_bF_buf12_bF_buf1_), .Y(_5322_) );
MUX2X1 MUX2X1_557 ( .gnd(gnd), .vdd(vdd), .A(_5322_), .B(_5317_), .S(_4036__bF_buf1), .Y(_5323_) );
MUX2X1 MUX2X1_558 ( .gnd(gnd), .vdd(vdd), .A(_5323_), .B(_5312_), .S(_4033__bF_buf3), .Y(_5324_) );
MUX2X1 MUX2X1_559 ( .gnd(gnd), .vdd(vdd), .A(_5324_), .B(_5301_), .S(raddr2_4_bF_buf2_), .Y(_5512__27_) );
NAND2X1 NAND2X1_1052 ( .gnd(gnd), .vdd(vdd), .A(regs_22__28_), .B(raddr2_0_bF_buf32_), .Y(_5325_) );
OAI21X1 OAI21X1_2046 ( .gnd(gnd), .vdd(vdd), .A(_1366_), .B(raddr2_0_bF_buf31_), .C(_5325_), .Y(_5326_) );
NAND2X1 NAND2X1_1053 ( .gnd(gnd), .vdd(vdd), .A(regs_20__28_), .B(raddr2_0_bF_buf30_), .Y(_5327_) );
OAI21X1 OAI21X1_2047 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(raddr2_0_bF_buf29_), .C(_5327_), .Y(_5328_) );
MUX2X1 MUX2X1_560 ( .gnd(gnd), .vdd(vdd), .A(_5328_), .B(_5326_), .S(raddr2_1_bF_buf11_), .Y(_5329_) );
NAND2X1 NAND2X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf0), .B(_5329_), .Y(_5330_) );
NAND2X1 NAND2X1_1055 ( .gnd(gnd), .vdd(vdd), .A(regs_18__28_), .B(raddr2_0_bF_buf28_), .Y(_5331_) );
OAI21X1 OAI21X1_2048 ( .gnd(gnd), .vdd(vdd), .A(_1563_), .B(raddr2_0_bF_buf27_), .C(_5331_), .Y(_5332_) );
NAND2X1 NAND2X1_1056 ( .gnd(gnd), .vdd(vdd), .A(regs_16__28_), .B(raddr2_0_bF_buf26_), .Y(_5333_) );
OAI21X1 OAI21X1_2049 ( .gnd(gnd), .vdd(vdd), .A(_1661_), .B(raddr2_0_bF_buf25_), .C(_5333_), .Y(_5334_) );
MUX2X1 MUX2X1_561 ( .gnd(gnd), .vdd(vdd), .A(_5334_), .B(_5332_), .S(raddr2_1_bF_buf10_), .Y(_5335_) );
AOI21X1 AOI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(raddr2_2_bF_buf3_), .B(_5335_), .C(_4033__bF_buf2), .Y(_5336_) );
OAI21X1 OAI21X1_2050 ( .gnd(gnd), .vdd(vdd), .A(_1199_), .B(raddr2_0_bF_buf24_), .C(raddr2_2_bF_buf2_), .Y(_5337_) );
AOI21X1 AOI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(regs_26__28_), .B(raddr2_0_bF_buf23_), .C(_5337_), .Y(_5338_) );
OAI21X1 OAI21X1_2051 ( .gnd(gnd), .vdd(vdd), .A(regs_30__28_), .B(raddr2_2_bF_buf1_), .C(_4038__bF_buf4), .Y(_5339_) );
OAI21X1 OAI21X1_2052 ( .gnd(gnd), .vdd(vdd), .A(_3843_), .B(raddr2_0_bF_buf22_), .C(raddr2_2_bF_buf0_), .Y(_5340_) );
AOI21X1 AOI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(regs_24__28_), .B(raddr2_0_bF_buf21_), .C(_5340_), .Y(_5341_) );
NOR2X1 NOR2X1_239 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf20_), .B(_3846_), .Y(_5342_) );
NAND2X1 NAND2X1_1057 ( .gnd(gnd), .vdd(vdd), .A(regs_28__28_), .B(raddr2_0_bF_buf19_), .Y(_5343_) );
NAND2X1 NAND2X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf8), .B(_5343_), .Y(_5344_) );
OAI21X1 OAI21X1_2053 ( .gnd(gnd), .vdd(vdd), .A(_5344_), .B(_5342_), .C(raddr2_1_bF_buf9_), .Y(_5345_) );
OAI22X1 OAI22X1_98 ( .gnd(gnd), .vdd(vdd), .A(_5338_), .B(_5339_), .C(_5345_), .D(_5341_), .Y(_5346_) );
AOI22X1 AOI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_5346_), .B(_4033__bF_buf1), .C(_5330_), .D(_5336_), .Y(_5347_) );
OAI21X1 OAI21X1_2054 ( .gnd(gnd), .vdd(vdd), .A(_3853_), .B(raddr2_0_bF_buf18_), .C(raddr2_1_bF_buf8_), .Y(_5348_) );
AOI21X1 AOI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(regs_4__28_), .B(raddr2_0_bF_buf17_), .C(_5348_), .Y(_5349_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(regs_6__28_), .B(raddr2_0_bF_buf16_), .Y(_5350_) );
OAI21X1 OAI21X1_2055 ( .gnd(gnd), .vdd(vdd), .A(_2157_), .B(raddr2_0_bF_buf15_), .C(_4038__bF_buf3), .Y(_5351_) );
OAI21X1 OAI21X1_2056 ( .gnd(gnd), .vdd(vdd), .A(_5351_), .B(_5350_), .C(_4036__bF_buf7), .Y(_5352_) );
OAI21X1 OAI21X1_2057 ( .gnd(gnd), .vdd(vdd), .A(_3859_), .B(raddr2_0_bF_buf14_), .C(raddr2_1_bF_buf7_), .Y(_5353_) );
AOI21X1 AOI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(regs_0__28_), .B(raddr2_0_bF_buf13_), .C(_5353_), .Y(_5354_) );
NOR2X1 NOR2X1_240 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf12_), .B(_3862_), .Y(_5355_) );
NAND2X1 NAND2X1_1059 ( .gnd(gnd), .vdd(vdd), .A(regs_2__28_), .B(raddr2_0_bF_buf11_), .Y(_5356_) );
NAND2X1 NAND2X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf2), .B(_5356_), .Y(_5357_) );
OAI21X1 OAI21X1_2058 ( .gnd(gnd), .vdd(vdd), .A(_5357_), .B(_5355_), .C(raddr2_2_bF_buf10_), .Y(_5358_) );
OAI22X1 OAI22X1_99 ( .gnd(gnd), .vdd(vdd), .A(_5354_), .B(_5358_), .C(_5352_), .D(_5349_), .Y(_5359_) );
NAND2X1 NAND2X1_1061 ( .gnd(gnd), .vdd(vdd), .A(regs_10__28_), .B(raddr2_0_bF_buf10_), .Y(_5360_) );
OAI21X1 OAI21X1_2059 ( .gnd(gnd), .vdd(vdd), .A(_1958_), .B(raddr2_0_bF_buf9_), .C(_5360_), .Y(_5361_) );
NAND2X1 NAND2X1_1062 ( .gnd(gnd), .vdd(vdd), .A(regs_8__28_), .B(raddr2_0_bF_buf8_), .Y(_5362_) );
OAI21X1 OAI21X1_2060 ( .gnd(gnd), .vdd(vdd), .A(_2056_), .B(raddr2_0_bF_buf7_), .C(_5362_), .Y(_5363_) );
MUX2X1 MUX2X1_562 ( .gnd(gnd), .vdd(vdd), .A(_5363_), .B(_5361_), .S(raddr2_1_bF_buf6_), .Y(_5364_) );
NAND2X1 NAND2X1_1063 ( .gnd(gnd), .vdd(vdd), .A(regs_14__28_), .B(raddr2_0_bF_buf6_), .Y(_5365_) );
OAI21X1 OAI21X1_2061 ( .gnd(gnd), .vdd(vdd), .A(_1761_), .B(raddr2_0_bF_buf5_), .C(_5365_), .Y(_5366_) );
NAND2X1 NAND2X1_1064 ( .gnd(gnd), .vdd(vdd), .A(regs_12__28_), .B(raddr2_0_bF_buf4_), .Y(_5367_) );
OAI21X1 OAI21X1_2062 ( .gnd(gnd), .vdd(vdd), .A(_1859_), .B(raddr2_0_bF_buf3_), .C(_5367_), .Y(_5368_) );
MUX2X1 MUX2X1_563 ( .gnd(gnd), .vdd(vdd), .A(_5368_), .B(_5366_), .S(raddr2_1_bF_buf5_), .Y(_5369_) );
MUX2X1 MUX2X1_564 ( .gnd(gnd), .vdd(vdd), .A(_5369_), .B(_5364_), .S(_4036__bF_buf6), .Y(_5370_) );
MUX2X1 MUX2X1_565 ( .gnd(gnd), .vdd(vdd), .A(_5370_), .B(_5359_), .S(_4033__bF_buf0), .Y(_5371_) );
MUX2X1 MUX2X1_566 ( .gnd(gnd), .vdd(vdd), .A(_5371_), .B(_5347_), .S(raddr2_4_bF_buf1_), .Y(_5512__28_) );
OAI21X1 OAI21X1_2063 ( .gnd(gnd), .vdd(vdd), .A(_3905_), .B(raddr2_0_bF_buf2_), .C(raddr2_1_bF_buf4_), .Y(_5372_) );
AOI21X1 AOI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(regs_4__29_), .B(raddr2_0_bF_buf1_), .C(_5372_), .Y(_5373_) );
AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(regs_6__29_), .B(raddr2_0_bF_buf0_), .Y(_5374_) );
OAI21X1 OAI21X1_2064 ( .gnd(gnd), .vdd(vdd), .A(_2159_), .B(raddr2_0_bF_buf96_), .C(_4038__bF_buf1), .Y(_5375_) );
OAI21X1 OAI21X1_2065 ( .gnd(gnd), .vdd(vdd), .A(_5375_), .B(_5374_), .C(_4036__bF_buf5), .Y(_5376_) );
OAI21X1 OAI21X1_2066 ( .gnd(gnd), .vdd(vdd), .A(_3911_), .B(raddr2_0_bF_buf95_), .C(raddr2_1_bF_buf3_), .Y(_5377_) );
AOI21X1 AOI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(regs_0__29_), .B(raddr2_0_bF_buf94_), .C(_5377_), .Y(_5378_) );
NOR2X1 NOR2X1_241 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf93_), .B(_3914_), .Y(_5379_) );
NAND2X1 NAND2X1_1065 ( .gnd(gnd), .vdd(vdd), .A(regs_2__29_), .B(raddr2_0_bF_buf92_), .Y(_5380_) );
NAND2X1 NAND2X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf0), .B(_5380_), .Y(_5381_) );
OAI21X1 OAI21X1_2067 ( .gnd(gnd), .vdd(vdd), .A(_5381_), .B(_5379_), .C(raddr2_2_bF_buf9_), .Y(_5382_) );
OAI22X1 OAI22X1_100 ( .gnd(gnd), .vdd(vdd), .A(_5378_), .B(_5382_), .C(_5376_), .D(_5373_), .Y(_5383_) );
NAND2X1 NAND2X1_1067 ( .gnd(gnd), .vdd(vdd), .A(regs_10__29_), .B(raddr2_0_bF_buf91_), .Y(_5384_) );
OAI21X1 OAI21X1_2068 ( .gnd(gnd), .vdd(vdd), .A(_1960_), .B(raddr2_0_bF_buf90_), .C(_5384_), .Y(_5385_) );
NAND2X1 NAND2X1_1068 ( .gnd(gnd), .vdd(vdd), .A(regs_8__29_), .B(raddr2_0_bF_buf89_), .Y(_5386_) );
OAI21X1 OAI21X1_2069 ( .gnd(gnd), .vdd(vdd), .A(_2058_), .B(raddr2_0_bF_buf88_), .C(_5386_), .Y(_5387_) );
MUX2X1 MUX2X1_567 ( .gnd(gnd), .vdd(vdd), .A(_5387_), .B(_5385_), .S(raddr2_1_bF_buf2_), .Y(_5388_) );
NAND2X1 NAND2X1_1069 ( .gnd(gnd), .vdd(vdd), .A(regs_14__29_), .B(raddr2_0_bF_buf87_), .Y(_5389_) );
OAI21X1 OAI21X1_2070 ( .gnd(gnd), .vdd(vdd), .A(_1763_), .B(raddr2_0_bF_buf86_), .C(_5389_), .Y(_5390_) );
NAND2X1 NAND2X1_1070 ( .gnd(gnd), .vdd(vdd), .A(regs_12__29_), .B(raddr2_0_bF_buf85_), .Y(_5391_) );
OAI21X1 OAI21X1_2071 ( .gnd(gnd), .vdd(vdd), .A(_1861_), .B(raddr2_0_bF_buf84_), .C(_5391_), .Y(_5392_) );
MUX2X1 MUX2X1_568 ( .gnd(gnd), .vdd(vdd), .A(_5392_), .B(_5390_), .S(raddr2_1_bF_buf1_), .Y(_5393_) );
MUX2X1 MUX2X1_569 ( .gnd(gnd), .vdd(vdd), .A(_5393_), .B(_5388_), .S(_4036__bF_buf4), .Y(_5394_) );
MUX2X1 MUX2X1_570 ( .gnd(gnd), .vdd(vdd), .A(_5394_), .B(_5383_), .S(_4033__bF_buf7), .Y(_5395_) );
OAI21X1 OAI21X1_2072 ( .gnd(gnd), .vdd(vdd), .A(_1663_), .B(raddr2_0_bF_buf83_), .C(raddr2_1_bF_buf0_), .Y(_5396_) );
AOI21X1 AOI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(regs_16__29_), .B(raddr2_0_bF_buf82_), .C(_5396_), .Y(_5397_) );
NOR2X1 NOR2X1_242 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf81_), .B(_1565_), .Y(_5398_) );
NAND2X1 NAND2X1_1071 ( .gnd(gnd), .vdd(vdd), .A(regs_18__29_), .B(raddr2_0_bF_buf80_), .Y(_5399_) );
NAND2X1 NAND2X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf8), .B(_5399_), .Y(_5400_) );
OAI21X1 OAI21X1_2073 ( .gnd(gnd), .vdd(vdd), .A(_5400_), .B(_5398_), .C(raddr2_2_bF_buf8_), .Y(_5401_) );
OAI21X1 OAI21X1_2074 ( .gnd(gnd), .vdd(vdd), .A(_1466_), .B(raddr2_0_bF_buf79_), .C(raddr2_1_bF_buf14_bF_buf0_), .Y(_5402_) );
AOI21X1 AOI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(regs_20__29_), .B(raddr2_0_bF_buf78_), .C(_5402_), .Y(_5403_) );
AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(regs_22__29_), .B(raddr2_0_bF_buf77_), .Y(_5404_) );
OAI21X1 OAI21X1_2075 ( .gnd(gnd), .vdd(vdd), .A(_1368_), .B(raddr2_0_bF_buf76_), .C(_4038__bF_buf7), .Y(_5405_) );
OAI21X1 OAI21X1_2076 ( .gnd(gnd), .vdd(vdd), .A(_5405_), .B(_5404_), .C(_4036__bF_buf3), .Y(_5406_) );
OAI22X1 OAI22X1_101 ( .gnd(gnd), .vdd(vdd), .A(_5397_), .B(_5401_), .C(_5406_), .D(_5403_), .Y(_5407_) );
NAND2X1 NAND2X1_1073 ( .gnd(gnd), .vdd(vdd), .A(regs_28__29_), .B(raddr2_0_bF_buf75_), .Y(_5408_) );
OAI21X1 OAI21X1_2077 ( .gnd(gnd), .vdd(vdd), .A(_3898_), .B(raddr2_0_bF_buf74_), .C(_5408_), .Y(_5409_) );
MUX2X1 MUX2X1_571 ( .gnd(gnd), .vdd(vdd), .A(_5409_), .B(regs_30__29_), .S(raddr2_1_bF_buf13_bF_buf0_), .Y(_5410_) );
NAND2X1 NAND2X1_1074 ( .gnd(gnd), .vdd(vdd), .A(regs_26__29_), .B(raddr2_0_bF_buf73_), .Y(_5411_) );
OAI21X1 OAI21X1_2078 ( .gnd(gnd), .vdd(vdd), .A(_1201_), .B(raddr2_0_bF_buf72_), .C(_5411_), .Y(_5412_) );
NAND2X1 NAND2X1_1075 ( .gnd(gnd), .vdd(vdd), .A(regs_24__29_), .B(raddr2_0_bF_buf71_), .Y(_5413_) );
OAI21X1 OAI21X1_2079 ( .gnd(gnd), .vdd(vdd), .A(_3895_), .B(raddr2_0_bF_buf70_), .C(_5413_), .Y(_5414_) );
MUX2X1 MUX2X1_572 ( .gnd(gnd), .vdd(vdd), .A(_5414_), .B(_5412_), .S(raddr2_1_bF_buf12_bF_buf0_), .Y(_5415_) );
MUX2X1 MUX2X1_573 ( .gnd(gnd), .vdd(vdd), .A(_5415_), .B(_5410_), .S(raddr2_2_bF_buf7_), .Y(_5416_) );
MUX2X1 MUX2X1_574 ( .gnd(gnd), .vdd(vdd), .A(_5416_), .B(_5407_), .S(_4033__bF_buf6), .Y(_5417_) );
MUX2X1 MUX2X1_575 ( .gnd(gnd), .vdd(vdd), .A(_5395_), .B(_5417_), .S(raddr2_4_bF_buf0_), .Y(_5512__29_) );
OAI21X1 OAI21X1_2080 ( .gnd(gnd), .vdd(vdd), .A(_3958_), .B(raddr2_0_bF_buf69_), .C(raddr2_1_bF_buf11_), .Y(_5418_) );
AOI21X1 AOI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(regs_4__30_), .B(raddr2_0_bF_buf68_), .C(_5418_), .Y(_5419_) );
AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(regs_6__30_), .B(raddr2_0_bF_buf67_), .Y(_5420_) );
OAI21X1 OAI21X1_2081 ( .gnd(gnd), .vdd(vdd), .A(_2161_), .B(raddr2_0_bF_buf66_), .C(_4038__bF_buf6), .Y(_5421_) );
OAI21X1 OAI21X1_2082 ( .gnd(gnd), .vdd(vdd), .A(_5421_), .B(_5420_), .C(_4036__bF_buf2), .Y(_5422_) );
OAI21X1 OAI21X1_2083 ( .gnd(gnd), .vdd(vdd), .A(_3965_), .B(raddr2_0_bF_buf65_), .C(raddr2_1_bF_buf10_), .Y(_5423_) );
AOI21X1 AOI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(regs_0__30_), .B(raddr2_0_bF_buf64_), .C(_5423_), .Y(_5424_) );
NOR2X1 NOR2X1_243 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf63_), .B(_3962_), .Y(_5425_) );
NAND2X1 NAND2X1_1076 ( .gnd(gnd), .vdd(vdd), .A(regs_2__30_), .B(raddr2_0_bF_buf62_), .Y(_5426_) );
NAND2X1 NAND2X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf5), .B(_5426_), .Y(_5427_) );
OAI21X1 OAI21X1_2084 ( .gnd(gnd), .vdd(vdd), .A(_5427_), .B(_5425_), .C(raddr2_2_bF_buf6_), .Y(_5428_) );
OAI22X1 OAI22X1_102 ( .gnd(gnd), .vdd(vdd), .A(_5424_), .B(_5428_), .C(_5422_), .D(_5419_), .Y(_5429_) );
NAND2X1 NAND2X1_1078 ( .gnd(gnd), .vdd(vdd), .A(regs_10__30_), .B(raddr2_0_bF_buf61_), .Y(_5430_) );
OAI21X1 OAI21X1_2085 ( .gnd(gnd), .vdd(vdd), .A(_1962_), .B(raddr2_0_bF_buf60_), .C(_5430_), .Y(_5431_) );
NAND2X1 NAND2X1_1079 ( .gnd(gnd), .vdd(vdd), .A(regs_8__30_), .B(raddr2_0_bF_buf59_), .Y(_5432_) );
OAI21X1 OAI21X1_2086 ( .gnd(gnd), .vdd(vdd), .A(_2060_), .B(raddr2_0_bF_buf58_), .C(_5432_), .Y(_5433_) );
MUX2X1 MUX2X1_576 ( .gnd(gnd), .vdd(vdd), .A(_5433_), .B(_5431_), .S(raddr2_1_bF_buf9_), .Y(_5434_) );
NAND2X1 NAND2X1_1080 ( .gnd(gnd), .vdd(vdd), .A(regs_14__30_), .B(raddr2_0_bF_buf57_), .Y(_5435_) );
OAI21X1 OAI21X1_2087 ( .gnd(gnd), .vdd(vdd), .A(_1765_), .B(raddr2_0_bF_buf56_), .C(_5435_), .Y(_5436_) );
NAND2X1 NAND2X1_1081 ( .gnd(gnd), .vdd(vdd), .A(regs_12__30_), .B(raddr2_0_bF_buf55_), .Y(_5437_) );
OAI21X1 OAI21X1_2088 ( .gnd(gnd), .vdd(vdd), .A(_1863_), .B(raddr2_0_bF_buf54_), .C(_5437_), .Y(_5438_) );
MUX2X1 MUX2X1_577 ( .gnd(gnd), .vdd(vdd), .A(_5438_), .B(_5436_), .S(raddr2_1_bF_buf8_), .Y(_5439_) );
MUX2X1 MUX2X1_578 ( .gnd(gnd), .vdd(vdd), .A(_5439_), .B(_5434_), .S(_4036__bF_buf1), .Y(_5440_) );
MUX2X1 MUX2X1_579 ( .gnd(gnd), .vdd(vdd), .A(_5440_), .B(_5429_), .S(_4033__bF_buf5), .Y(_5441_) );
OAI21X1 OAI21X1_2089 ( .gnd(gnd), .vdd(vdd), .A(_1665_), .B(raddr2_0_bF_buf53_), .C(raddr2_1_bF_buf7_), .Y(_5442_) );
AOI21X1 AOI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(regs_16__30_), .B(raddr2_0_bF_buf52_), .C(_5442_), .Y(_5443_) );
NOR2X1 NOR2X1_244 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf51_), .B(_1567_), .Y(_5444_) );
NAND2X1 NAND2X1_1082 ( .gnd(gnd), .vdd(vdd), .A(regs_18__30_), .B(raddr2_0_bF_buf50_), .Y(_5445_) );
NAND2X1 NAND2X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf4), .B(_5445_), .Y(_5446_) );
OAI21X1 OAI21X1_2090 ( .gnd(gnd), .vdd(vdd), .A(_5446_), .B(_5444_), .C(raddr2_2_bF_buf5_), .Y(_5447_) );
OAI21X1 OAI21X1_2091 ( .gnd(gnd), .vdd(vdd), .A(_1468_), .B(raddr2_0_bF_buf49_), .C(raddr2_1_bF_buf6_), .Y(_5448_) );
AOI21X1 AOI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(regs_20__30_), .B(raddr2_0_bF_buf48_), .C(_5448_), .Y(_5449_) );
AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(regs_22__30_), .B(raddr2_0_bF_buf47_), .Y(_5450_) );
OAI21X1 OAI21X1_2092 ( .gnd(gnd), .vdd(vdd), .A(_1370_), .B(raddr2_0_bF_buf46_), .C(_4038__bF_buf3), .Y(_5451_) );
OAI21X1 OAI21X1_2093 ( .gnd(gnd), .vdd(vdd), .A(_5451_), .B(_5450_), .C(_4036__bF_buf0), .Y(_5452_) );
OAI22X1 OAI22X1_103 ( .gnd(gnd), .vdd(vdd), .A(_5443_), .B(_5447_), .C(_5452_), .D(_5449_), .Y(_5453_) );
NAND2X1 NAND2X1_1084 ( .gnd(gnd), .vdd(vdd), .A(regs_28__30_), .B(raddr2_0_bF_buf45_), .Y(_5454_) );
OAI21X1 OAI21X1_2094 ( .gnd(gnd), .vdd(vdd), .A(_3944_), .B(raddr2_0_bF_buf44_), .C(_5454_), .Y(_5455_) );
MUX2X1 MUX2X1_580 ( .gnd(gnd), .vdd(vdd), .A(_5455_), .B(regs_30__30_), .S(raddr2_1_bF_buf5_), .Y(_5456_) );
NAND2X1 NAND2X1_1085 ( .gnd(gnd), .vdd(vdd), .A(regs_26__30_), .B(raddr2_0_bF_buf43_), .Y(_5457_) );
OAI21X1 OAI21X1_2095 ( .gnd(gnd), .vdd(vdd), .A(_1203_), .B(raddr2_0_bF_buf42_), .C(_5457_), .Y(_5458_) );
NAND2X1 NAND2X1_1086 ( .gnd(gnd), .vdd(vdd), .A(regs_24__30_), .B(raddr2_0_bF_buf41_), .Y(_5459_) );
OAI21X1 OAI21X1_2096 ( .gnd(gnd), .vdd(vdd), .A(_3950_), .B(raddr2_0_bF_buf40_), .C(_5459_), .Y(_5460_) );
MUX2X1 MUX2X1_581 ( .gnd(gnd), .vdd(vdd), .A(_5460_), .B(_5458_), .S(raddr2_1_bF_buf4_), .Y(_5461_) );
MUX2X1 MUX2X1_582 ( .gnd(gnd), .vdd(vdd), .A(_5461_), .B(_5456_), .S(raddr2_2_bF_buf4_), .Y(_5462_) );
MUX2X1 MUX2X1_583 ( .gnd(gnd), .vdd(vdd), .A(_5462_), .B(_5453_), .S(_4033__bF_buf4), .Y(_5463_) );
MUX2X1 MUX2X1_584 ( .gnd(gnd), .vdd(vdd), .A(_5441_), .B(_5463_), .S(raddr2_4_bF_buf4_), .Y(_5512__30_) );
NAND2X1 NAND2X1_1087 ( .gnd(gnd), .vdd(vdd), .A(regs_22__31_), .B(raddr2_0_bF_buf39_), .Y(_5464_) );
OAI21X1 OAI21X1_2097 ( .gnd(gnd), .vdd(vdd), .A(_1372_), .B(raddr2_0_bF_buf38_), .C(_5464_), .Y(_5465_) );
NAND2X1 NAND2X1_1088 ( .gnd(gnd), .vdd(vdd), .A(regs_20__31_), .B(raddr2_0_bF_buf37_), .Y(_5466_) );
OAI21X1 OAI21X1_2098 ( .gnd(gnd), .vdd(vdd), .A(_1470_), .B(raddr2_0_bF_buf36_), .C(_5466_), .Y(_5467_) );
MUX2X1 MUX2X1_585 ( .gnd(gnd), .vdd(vdd), .A(_5467_), .B(_5465_), .S(raddr2_1_bF_buf3_), .Y(_5468_) );
NAND2X1 NAND2X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf8), .B(_5468_), .Y(_5469_) );
NAND2X1 NAND2X1_1090 ( .gnd(gnd), .vdd(vdd), .A(regs_18__31_), .B(raddr2_0_bF_buf35_), .Y(_5470_) );
OAI21X1 OAI21X1_2099 ( .gnd(gnd), .vdd(vdd), .A(_1569_), .B(raddr2_0_bF_buf34_), .C(_5470_), .Y(_5471_) );
NAND2X1 NAND2X1_1091 ( .gnd(gnd), .vdd(vdd), .A(regs_16__31_), .B(raddr2_0_bF_buf33_), .Y(_5472_) );
OAI21X1 OAI21X1_2100 ( .gnd(gnd), .vdd(vdd), .A(_1667_), .B(raddr2_0_bF_buf32_), .C(_5472_), .Y(_5473_) );
MUX2X1 MUX2X1_586 ( .gnd(gnd), .vdd(vdd), .A(_5473_), .B(_5471_), .S(raddr2_1_bF_buf2_), .Y(_5474_) );
AOI21X1 AOI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(raddr2_2_bF_buf3_), .B(_5474_), .C(_4033__bF_buf3), .Y(_5475_) );
OAI21X1 OAI21X1_2101 ( .gnd(gnd), .vdd(vdd), .A(_1205_), .B(raddr2_0_bF_buf31_), .C(raddr2_2_bF_buf2_), .Y(_5476_) );
AOI21X1 AOI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(regs_26__31_), .B(raddr2_0_bF_buf30_), .C(_5476_), .Y(_5477_) );
OAI21X1 OAI21X1_2102 ( .gnd(gnd), .vdd(vdd), .A(regs_30__31_), .B(raddr2_2_bF_buf1_), .C(_4038__bF_buf2), .Y(_5478_) );
OAI21X1 OAI21X1_2103 ( .gnd(gnd), .vdd(vdd), .A(_4027_), .B(raddr2_0_bF_buf29_), .C(raddr2_2_bF_buf0_), .Y(_5479_) );
AOI21X1 AOI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(regs_24__31_), .B(raddr2_0_bF_buf28_), .C(_5479_), .Y(_5480_) );
NOR2X1 NOR2X1_245 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf27_), .B(_4021_), .Y(_5481_) );
NAND2X1 NAND2X1_1092 ( .gnd(gnd), .vdd(vdd), .A(regs_28__31_), .B(raddr2_0_bF_buf26_), .Y(_5482_) );
NAND2X1 NAND2X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_4036__bF_buf7), .B(_5482_), .Y(_5483_) );
OAI21X1 OAI21X1_2104 ( .gnd(gnd), .vdd(vdd), .A(_5483_), .B(_5481_), .C(raddr2_1_bF_buf1_), .Y(_5484_) );
OAI22X1 OAI22X1_104 ( .gnd(gnd), .vdd(vdd), .A(_5477_), .B(_5478_), .C(_5484_), .D(_5480_), .Y(_5485_) );
AOI22X1 AOI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_5485_), .B(_4033__bF_buf2), .C(_5469_), .D(_5475_), .Y(_5486_) );
OAI21X1 OAI21X1_2105 ( .gnd(gnd), .vdd(vdd), .A(_3982_), .B(raddr2_0_bF_buf25_), .C(raddr2_1_bF_buf0_), .Y(_5487_) );
AOI21X1 AOI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(regs_4__31_), .B(raddr2_0_bF_buf24_), .C(_5487_), .Y(_5488_) );
AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(regs_6__31_), .B(raddr2_0_bF_buf23_), .Y(_5489_) );
OAI21X1 OAI21X1_2106 ( .gnd(gnd), .vdd(vdd), .A(_2163_), .B(raddr2_0_bF_buf22_), .C(_4038__bF_buf1), .Y(_5490_) );
OAI21X1 OAI21X1_2107 ( .gnd(gnd), .vdd(vdd), .A(_5490_), .B(_5489_), .C(_4036__bF_buf6), .Y(_5491_) );
OAI21X1 OAI21X1_2108 ( .gnd(gnd), .vdd(vdd), .A(_3988_), .B(raddr2_0_bF_buf21_), .C(raddr2_1_bF_buf14_bF_buf3_), .Y(_5492_) );
AOI21X1 AOI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(regs_0__31_), .B(raddr2_0_bF_buf20_), .C(_5492_), .Y(_5493_) );
NOR2X1 NOR2X1_246 ( .gnd(gnd), .vdd(vdd), .A(raddr2_0_bF_buf19_), .B(_3991_), .Y(_5494_) );
NAND2X1 NAND2X1_1094 ( .gnd(gnd), .vdd(vdd), .A(regs_2__31_), .B(raddr2_0_bF_buf18_), .Y(_5495_) );
NAND2X1 NAND2X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_4038__bF_buf0), .B(_5495_), .Y(_5496_) );
OAI21X1 OAI21X1_2109 ( .gnd(gnd), .vdd(vdd), .A(_5496_), .B(_5494_), .C(raddr2_2_bF_buf10_), .Y(_5497_) );
OAI22X1 OAI22X1_105 ( .gnd(gnd), .vdd(vdd), .A(_5493_), .B(_5497_), .C(_5491_), .D(_5488_), .Y(_5498_) );
NAND2X1 NAND2X1_1096 ( .gnd(gnd), .vdd(vdd), .A(regs_10__31_), .B(raddr2_0_bF_buf17_), .Y(_5499_) );
OAI21X1 OAI21X1_2110 ( .gnd(gnd), .vdd(vdd), .A(_1964_), .B(raddr2_0_bF_buf16_), .C(_5499_), .Y(_5500_) );
NAND2X1 NAND2X1_1097 ( .gnd(gnd), .vdd(vdd), .A(regs_8__31_), .B(raddr2_0_bF_buf15_), .Y(_5501_) );
OAI21X1 OAI21X1_2111 ( .gnd(gnd), .vdd(vdd), .A(_2062_), .B(raddr2_0_bF_buf14_), .C(_5501_), .Y(_5502_) );
MUX2X1 MUX2X1_587 ( .gnd(gnd), .vdd(vdd), .A(_5502_), .B(_5500_), .S(raddr2_1_bF_buf13_bF_buf3_), .Y(_5503_) );
NAND2X1 NAND2X1_1098 ( .gnd(gnd), .vdd(vdd), .A(regs_14__31_), .B(raddr2_0_bF_buf13_), .Y(_5504_) );
OAI21X1 OAI21X1_2112 ( .gnd(gnd), .vdd(vdd), .A(_1767_), .B(raddr2_0_bF_buf12_), .C(_5504_), .Y(_5505_) );
NAND2X1 NAND2X1_1099 ( .gnd(gnd), .vdd(vdd), .A(regs_12__31_), .B(raddr2_0_bF_buf11_), .Y(_5506_) );
OAI21X1 OAI21X1_2113 ( .gnd(gnd), .vdd(vdd), .A(_1865_), .B(raddr2_0_bF_buf10_), .C(_5506_), .Y(_5507_) );
MUX2X1 MUX2X1_588 ( .gnd(gnd), .vdd(vdd), .A(_5507_), .B(_5505_), .S(raddr2_1_bF_buf12_bF_buf3_), .Y(_5508_) );
MUX2X1 MUX2X1_589 ( .gnd(gnd), .vdd(vdd), .A(_5508_), .B(_5503_), .S(_4036__bF_buf5), .Y(_5509_) );
MUX2X1 MUX2X1_590 ( .gnd(gnd), .vdd(vdd), .A(_5509_), .B(_5498_), .S(_4033__bF_buf1), .Y(_5510_) );
MUX2X1 MUX2X1_591 ( .gnd(gnd), .vdd(vdd), .A(_5510_), .B(_5486_), .S(raddr2_4_bF_buf3_), .Y(_5512__31_) );
INVX8 INVX8_8 ( .gnd(gnd), .vdd(vdd), .A(wdata[0]), .Y(_992_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(waddr[4]), .Y(_993_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(waddr[3]), .Y(_994_) );
NAND2X1 NAND2X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_993_), .B(_994_), .Y(_995_) );
NOR2X1 NOR2X1_247 ( .gnd(gnd), .vdd(vdd), .A(waddr[2]), .B(_995_), .Y(_996_) );
NAND2X1 NAND2X1_1101 ( .gnd(gnd), .vdd(vdd), .A(waddr[0]), .B(wen), .Y(_997_) );
NOR2X1 NOR2X1_248 ( .gnd(gnd), .vdd(vdd), .A(waddr[1]), .B(_997_), .Y(_998_) );
NAND2X1 NAND2X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_998_), .B(_996_), .Y(_999_) );
INVX8 INVX8_9 ( .gnd(gnd), .vdd(vdd), .A(_996_), .Y(_1000_) );
INVX8 INVX8_10 ( .gnd(gnd), .vdd(vdd), .A(_998_), .Y(_1001_) );
OAI21X1 OAI21X1_2114 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf7), .B(_1001__bF_buf1), .C(regs_30__0_), .Y(_1002_) );
OAI21X1 OAI21X1_2115 ( .gnd(gnd), .vdd(vdd), .A(_992__bF_buf0), .B(_999__bF_buf4), .C(_1002_), .Y(_736_) );
INVX8 INVX8_11 ( .gnd(gnd), .vdd(vdd), .A(wdata[1]), .Y(_1003_) );
OAI21X1 OAI21X1_2116 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf6), .B(_1001__bF_buf0), .C(regs_30__1_), .Y(_1004_) );
OAI21X1 OAI21X1_2117 ( .gnd(gnd), .vdd(vdd), .A(_1003__bF_buf0), .B(_999__bF_buf3), .C(_1004_), .Y(_747_) );
INVX8 INVX8_12 ( .gnd(gnd), .vdd(vdd), .A(wdata[2]), .Y(_1005_) );
OAI21X1 OAI21X1_2118 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf5), .B(_1001__bF_buf9), .C(regs_30__2_), .Y(_1006_) );
OAI21X1 OAI21X1_2119 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf0), .B(_999__bF_buf2), .C(_1006_), .Y(_758_) );
INVX8 INVX8_13 ( .gnd(gnd), .vdd(vdd), .A(wdata[3]), .Y(_1007_) );
OAI21X1 OAI21X1_2120 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_1001__bF_buf8), .C(regs_30__3_), .Y(_1008_) );
OAI21X1 OAI21X1_2121 ( .gnd(gnd), .vdd(vdd), .A(_1007__bF_buf0), .B(_999__bF_buf1), .C(_1008_), .Y(_761_) );
INVX8 INVX8_14 ( .gnd(gnd), .vdd(vdd), .A(wdata[4]), .Y(_1009_) );
OAI21X1 OAI21X1_2122 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf3), .B(_1001__bF_buf7), .C(regs_30__4_), .Y(_1010_) );
OAI21X1 OAI21X1_2123 ( .gnd(gnd), .vdd(vdd), .A(_1009__bF_buf3), .B(_999__bF_buf0), .C(_1010_), .Y(_762_) );
INVX8 INVX8_15 ( .gnd(gnd), .vdd(vdd), .A(wdata[5]), .Y(_1011_) );
OAI21X1 OAI21X1_2124 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf2), .B(_1001__bF_buf6), .C(regs_30__5_), .Y(_1012_) );
OAI21X1 OAI21X1_2125 ( .gnd(gnd), .vdd(vdd), .A(_1011__bF_buf3), .B(_999__bF_buf4), .C(_1012_), .Y(_763_) );
INVX8 INVX8_16 ( .gnd(gnd), .vdd(vdd), .A(wdata[6]), .Y(_1013_) );
OAI21X1 OAI21X1_2126 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1001__bF_buf5), .C(regs_30__6_), .Y(_1014_) );
OAI21X1 OAI21X1_2127 ( .gnd(gnd), .vdd(vdd), .A(_1013__bF_buf3), .B(_999__bF_buf3), .C(_1014_), .Y(_764_) );
INVX8 INVX8_17 ( .gnd(gnd), .vdd(vdd), .A(wdata[7]), .Y(_1015_) );
OAI21X1 OAI21X1_2128 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf0), .B(_1001__bF_buf4), .C(regs_30__7_), .Y(_1016_) );
OAI21X1 OAI21X1_2129 ( .gnd(gnd), .vdd(vdd), .A(_1015__bF_buf3), .B(_999__bF_buf2), .C(_1016_), .Y(_765_) );
INVX8 INVX8_18 ( .gnd(gnd), .vdd(vdd), .A(wdata[8]), .Y(_1017_) );
OAI21X1 OAI21X1_2130 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf7), .B(_1001__bF_buf3), .C(regs_30__8_), .Y(_1018_) );
OAI21X1 OAI21X1_2131 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf3), .B(_999__bF_buf1), .C(_1018_), .Y(_766_) );
INVX8 INVX8_19 ( .gnd(gnd), .vdd(vdd), .A(wdata[9]), .Y(_1019_) );
OAI21X1 OAI21X1_2132 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf6), .B(_1001__bF_buf2), .C(regs_30__9_), .Y(_1020_) );
OAI21X1 OAI21X1_2133 ( .gnd(gnd), .vdd(vdd), .A(_1019__bF_buf3), .B(_999__bF_buf0), .C(_1020_), .Y(_767_) );
INVX8 INVX8_20 ( .gnd(gnd), .vdd(vdd), .A(wdata[10]), .Y(_1021_) );
OAI21X1 OAI21X1_2134 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf5), .B(_1001__bF_buf1), .C(regs_30__10_), .Y(_1022_) );
OAI21X1 OAI21X1_2135 ( .gnd(gnd), .vdd(vdd), .A(_1021__bF_buf3), .B(_999__bF_buf4), .C(_1022_), .Y(_737_) );
INVX8 INVX8_21 ( .gnd(gnd), .vdd(vdd), .A(wdata[11]), .Y(_1023_) );
OAI21X1 OAI21X1_2136 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_1001__bF_buf0), .C(regs_30__11_), .Y(_1024_) );
OAI21X1 OAI21X1_2137 ( .gnd(gnd), .vdd(vdd), .A(_1023__bF_buf3), .B(_999__bF_buf3), .C(_1024_), .Y(_738_) );
INVX8 INVX8_22 ( .gnd(gnd), .vdd(vdd), .A(wdata[12]), .Y(_1025_) );
OAI21X1 OAI21X1_2138 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf3), .B(_1001__bF_buf9), .C(regs_30__12_), .Y(_1026_) );
OAI21X1 OAI21X1_2139 ( .gnd(gnd), .vdd(vdd), .A(_1025__bF_buf3), .B(_999__bF_buf2), .C(_1026_), .Y(_739_) );
INVX8 INVX8_23 ( .gnd(gnd), .vdd(vdd), .A(wdata[13]), .Y(_1027_) );
OAI21X1 OAI21X1_2140 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf2), .B(_1001__bF_buf8), .C(regs_30__13_), .Y(_1028_) );
OAI21X1 OAI21X1_2141 ( .gnd(gnd), .vdd(vdd), .A(_1027__bF_buf3), .B(_999__bF_buf1), .C(_1028_), .Y(_740_) );
INVX8 INVX8_24 ( .gnd(gnd), .vdd(vdd), .A(wdata[14]), .Y(_1029_) );
OAI21X1 OAI21X1_2142 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1001__bF_buf7), .C(regs_30__14_), .Y(_1030_) );
OAI21X1 OAI21X1_2143 ( .gnd(gnd), .vdd(vdd), .A(_1029__bF_buf3), .B(_999__bF_buf0), .C(_1030_), .Y(_741_) );
INVX8 INVX8_25 ( .gnd(gnd), .vdd(vdd), .A(wdata[15]), .Y(_1031_) );
OAI21X1 OAI21X1_2144 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf0), .B(_1001__bF_buf6), .C(regs_30__15_), .Y(_1032_) );
OAI21X1 OAI21X1_2145 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf3), .B(_999__bF_buf4), .C(_1032_), .Y(_742_) );
INVX8 INVX8_26 ( .gnd(gnd), .vdd(vdd), .A(wdata[16]), .Y(_1033_) );
OAI21X1 OAI21X1_2146 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf7), .B(_1001__bF_buf5), .C(regs_30__16_), .Y(_1034_) );
OAI21X1 OAI21X1_2147 ( .gnd(gnd), .vdd(vdd), .A(_1033__bF_buf3), .B(_999__bF_buf3), .C(_1034_), .Y(_743_) );
INVX8 INVX8_27 ( .gnd(gnd), .vdd(vdd), .A(wdata[17]), .Y(_1035_) );
OAI21X1 OAI21X1_2148 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf6), .B(_1001__bF_buf4), .C(regs_30__17_), .Y(_1036_) );
OAI21X1 OAI21X1_2149 ( .gnd(gnd), .vdd(vdd), .A(_1035__bF_buf3), .B(_999__bF_buf2), .C(_1036_), .Y(_744_) );
INVX8 INVX8_28 ( .gnd(gnd), .vdd(vdd), .A(wdata[18]), .Y(_1037_) );
OAI21X1 OAI21X1_2150 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf5), .B(_1001__bF_buf3), .C(regs_30__18_), .Y(_1038_) );
OAI21X1 OAI21X1_2151 ( .gnd(gnd), .vdd(vdd), .A(_1037__bF_buf3), .B(_999__bF_buf1), .C(_1038_), .Y(_745_) );
INVX8 INVX8_29 ( .gnd(gnd), .vdd(vdd), .A(wdata[19]), .Y(_1039_) );
OAI21X1 OAI21X1_2152 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_1001__bF_buf2), .C(regs_30__19_), .Y(_1040_) );
OAI21X1 OAI21X1_2153 ( .gnd(gnd), .vdd(vdd), .A(_1039__bF_buf3), .B(_999__bF_buf0), .C(_1040_), .Y(_746_) );
INVX8 INVX8_30 ( .gnd(gnd), .vdd(vdd), .A(wdata[20]), .Y(_1041_) );
OAI21X1 OAI21X1_2154 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf3), .B(_1001__bF_buf1), .C(regs_30__20_), .Y(_1042_) );
OAI21X1 OAI21X1_2155 ( .gnd(gnd), .vdd(vdd), .A(_1041__bF_buf3), .B(_999__bF_buf4), .C(_1042_), .Y(_748_) );
INVX8 INVX8_31 ( .gnd(gnd), .vdd(vdd), .A(wdata[21]), .Y(_1043_) );
OAI21X1 OAI21X1_2156 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf2), .B(_1001__bF_buf0), .C(regs_30__21_), .Y(_1044_) );
OAI21X1 OAI21X1_2157 ( .gnd(gnd), .vdd(vdd), .A(_1043__bF_buf3), .B(_999__bF_buf3), .C(_1044_), .Y(_749_) );
INVX8 INVX8_32 ( .gnd(gnd), .vdd(vdd), .A(wdata[22]), .Y(_1045_) );
OAI21X1 OAI21X1_2158 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1001__bF_buf9), .C(regs_30__22_), .Y(_1046_) );
OAI21X1 OAI21X1_2159 ( .gnd(gnd), .vdd(vdd), .A(_1045__bF_buf3), .B(_999__bF_buf2), .C(_1046_), .Y(_750_) );
INVX8 INVX8_33 ( .gnd(gnd), .vdd(vdd), .A(wdata[23]), .Y(_1047_) );
OAI21X1 OAI21X1_2160 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf0), .B(_1001__bF_buf8), .C(regs_30__23_), .Y(_1048_) );
OAI21X1 OAI21X1_2161 ( .gnd(gnd), .vdd(vdd), .A(_1047__bF_buf3), .B(_999__bF_buf1), .C(_1048_), .Y(_751_) );
INVX8 INVX8_34 ( .gnd(gnd), .vdd(vdd), .A(wdata[24]), .Y(_1049_) );
OAI21X1 OAI21X1_2162 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf7), .B(_1001__bF_buf7), .C(regs_30__24_), .Y(_1050_) );
OAI21X1 OAI21X1_2163 ( .gnd(gnd), .vdd(vdd), .A(_1049__bF_buf3), .B(_999__bF_buf0), .C(_1050_), .Y(_752_) );
INVX8 INVX8_35 ( .gnd(gnd), .vdd(vdd), .A(wdata[25]), .Y(_1051_) );
OAI21X1 OAI21X1_2164 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf6), .B(_1001__bF_buf6), .C(regs_30__25_), .Y(_1052_) );
OAI21X1 OAI21X1_2165 ( .gnd(gnd), .vdd(vdd), .A(_1051__bF_buf3), .B(_999__bF_buf4), .C(_1052_), .Y(_753_) );
INVX8 INVX8_36 ( .gnd(gnd), .vdd(vdd), .A(wdata[26]), .Y(_1053_) );
OAI21X1 OAI21X1_2166 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf5), .B(_1001__bF_buf5), .C(regs_30__26_), .Y(_1054_) );
OAI21X1 OAI21X1_2167 ( .gnd(gnd), .vdd(vdd), .A(_1053__bF_buf3), .B(_999__bF_buf3), .C(_1054_), .Y(_754_) );
INVX8 INVX8_37 ( .gnd(gnd), .vdd(vdd), .A(wdata[27]), .Y(_1055_) );
OAI21X1 OAI21X1_2168 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_1001__bF_buf4), .C(regs_30__27_), .Y(_1056_) );
OAI21X1 OAI21X1_2169 ( .gnd(gnd), .vdd(vdd), .A(_1055__bF_buf3), .B(_999__bF_buf2), .C(_1056_), .Y(_755_) );
INVX8 INVX8_38 ( .gnd(gnd), .vdd(vdd), .A(wdata[28]), .Y(_1057_) );
OAI21X1 OAI21X1_2170 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf3), .B(_1001__bF_buf3), .C(regs_30__28_), .Y(_1058_) );
OAI21X1 OAI21X1_2171 ( .gnd(gnd), .vdd(vdd), .A(_1057__bF_buf3), .B(_999__bF_buf1), .C(_1058_), .Y(_756_) );
INVX8 INVX8_39 ( .gnd(gnd), .vdd(vdd), .A(wdata[29]), .Y(_1059_) );
OAI21X1 OAI21X1_2172 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf2), .B(_1001__bF_buf2), .C(regs_30__29_), .Y(_1060_) );
OAI21X1 OAI21X1_2173 ( .gnd(gnd), .vdd(vdd), .A(_1059__bF_buf3), .B(_999__bF_buf0), .C(_1060_), .Y(_757_) );
INVX8 INVX8_40 ( .gnd(gnd), .vdd(vdd), .A(wdata[30]), .Y(_1061_) );
OAI21X1 OAI21X1_2174 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1001__bF_buf1), .C(regs_30__30_), .Y(_1062_) );
OAI21X1 OAI21X1_2175 ( .gnd(gnd), .vdd(vdd), .A(_1061__bF_buf3), .B(_999__bF_buf4), .C(_1062_), .Y(_759_) );
INVX8 INVX8_41 ( .gnd(gnd), .vdd(vdd), .A(wdata[31]), .Y(_1063_) );
OAI21X1 OAI21X1_2176 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf0), .B(_1001__bF_buf0), .C(regs_30__31_), .Y(_1064_) );
OAI21X1 OAI21X1_2177 ( .gnd(gnd), .vdd(vdd), .A(_1063__bF_buf3), .B(_999__bF_buf3), .C(_1064_), .Y(_760_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(wen), .Y(_1065_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(waddr[0]), .Y(_1066_) );
NAND2X1 NAND2X1_1103 ( .gnd(gnd), .vdd(vdd), .A(waddr[1]), .B(_1066_), .Y(_1067_) );
NOR2X1 NOR2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1065_), .B(_1067_), .Y(_1068_) );
NAND2X1 NAND2X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_996_), .Y(_1069_) );
INVX8 INVX8_42 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .Y(_1070_) );
OAI21X1 OAI21X1_2178 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf7), .B(_1070__bF_buf8), .C(regs_29__0_), .Y(_1071_) );
OAI21X1 OAI21X1_2179 ( .gnd(gnd), .vdd(vdd), .A(_992__bF_buf3), .B(_1069__bF_buf4), .C(_1071_), .Y(_672_) );
OAI21X1 OAI21X1_2180 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf6), .B(_1070__bF_buf7), .C(regs_29__1_), .Y(_1072_) );
OAI21X1 OAI21X1_2181 ( .gnd(gnd), .vdd(vdd), .A(_1003__bF_buf3), .B(_1069__bF_buf3), .C(_1072_), .Y(_683_) );
OAI21X1 OAI21X1_2182 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf5), .B(_1070__bF_buf6), .C(regs_29__2_), .Y(_1073_) );
OAI21X1 OAI21X1_2183 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf3), .B(_1069__bF_buf2), .C(_1073_), .Y(_694_) );
OAI21X1 OAI21X1_2184 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_1070__bF_buf5), .C(regs_29__3_), .Y(_1074_) );
OAI21X1 OAI21X1_2185 ( .gnd(gnd), .vdd(vdd), .A(_1007__bF_buf3), .B(_1069__bF_buf1), .C(_1074_), .Y(_697_) );
OAI21X1 OAI21X1_2186 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf3), .B(_1070__bF_buf4), .C(regs_29__4_), .Y(_1075_) );
OAI21X1 OAI21X1_2187 ( .gnd(gnd), .vdd(vdd), .A(_1009__bF_buf2), .B(_1069__bF_buf0), .C(_1075_), .Y(_698_) );
OAI21X1 OAI21X1_2188 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf2), .B(_1070__bF_buf3), .C(regs_29__5_), .Y(_1076_) );
OAI21X1 OAI21X1_2189 ( .gnd(gnd), .vdd(vdd), .A(_1011__bF_buf2), .B(_1069__bF_buf4), .C(_1076_), .Y(_699_) );
OAI21X1 OAI21X1_2190 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1070__bF_buf2), .C(regs_29__6_), .Y(_1077_) );
OAI21X1 OAI21X1_2191 ( .gnd(gnd), .vdd(vdd), .A(_1013__bF_buf2), .B(_1069__bF_buf3), .C(_1077_), .Y(_700_) );
OAI21X1 OAI21X1_2192 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf0), .B(_1070__bF_buf1), .C(regs_29__7_), .Y(_1078_) );
OAI21X1 OAI21X1_2193 ( .gnd(gnd), .vdd(vdd), .A(_1015__bF_buf2), .B(_1069__bF_buf2), .C(_1078_), .Y(_701_) );
OAI21X1 OAI21X1_2194 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf7), .B(_1070__bF_buf0), .C(regs_29__8_), .Y(_1079_) );
OAI21X1 OAI21X1_2195 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf2), .B(_1069__bF_buf1), .C(_1079_), .Y(_702_) );
OAI21X1 OAI21X1_2196 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf6), .B(_1070__bF_buf10), .C(regs_29__9_), .Y(_1080_) );
OAI21X1 OAI21X1_2197 ( .gnd(gnd), .vdd(vdd), .A(_1019__bF_buf2), .B(_1069__bF_buf0), .C(_1080_), .Y(_703_) );
OAI21X1 OAI21X1_2198 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf5), .B(_1070__bF_buf9), .C(regs_29__10_), .Y(_1081_) );
OAI21X1 OAI21X1_2199 ( .gnd(gnd), .vdd(vdd), .A(_1021__bF_buf2), .B(_1069__bF_buf4), .C(_1081_), .Y(_673_) );
OAI21X1 OAI21X1_2200 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_1070__bF_buf8), .C(regs_29__11_), .Y(_1082_) );
OAI21X1 OAI21X1_2201 ( .gnd(gnd), .vdd(vdd), .A(_1023__bF_buf2), .B(_1069__bF_buf3), .C(_1082_), .Y(_674_) );
OAI21X1 OAI21X1_2202 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf3), .B(_1070__bF_buf7), .C(regs_29__12_), .Y(_1083_) );
OAI21X1 OAI21X1_2203 ( .gnd(gnd), .vdd(vdd), .A(_1025__bF_buf2), .B(_1069__bF_buf2), .C(_1083_), .Y(_675_) );
OAI21X1 OAI21X1_2204 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf2), .B(_1070__bF_buf6), .C(regs_29__13_), .Y(_1084_) );
OAI21X1 OAI21X1_2205 ( .gnd(gnd), .vdd(vdd), .A(_1027__bF_buf2), .B(_1069__bF_buf1), .C(_1084_), .Y(_676_) );
OAI21X1 OAI21X1_2206 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1070__bF_buf5), .C(regs_29__14_), .Y(_1085_) );
OAI21X1 OAI21X1_2207 ( .gnd(gnd), .vdd(vdd), .A(_1029__bF_buf2), .B(_1069__bF_buf0), .C(_1085_), .Y(_677_) );
OAI21X1 OAI21X1_2208 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf0), .B(_1070__bF_buf4), .C(regs_29__15_), .Y(_1086_) );
OAI21X1 OAI21X1_2209 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf2), .B(_1069__bF_buf4), .C(_1086_), .Y(_678_) );
OAI21X1 OAI21X1_2210 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf7), .B(_1070__bF_buf3), .C(regs_29__16_), .Y(_1087_) );
OAI21X1 OAI21X1_2211 ( .gnd(gnd), .vdd(vdd), .A(_1033__bF_buf2), .B(_1069__bF_buf3), .C(_1087_), .Y(_679_) );
OAI21X1 OAI21X1_2212 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf6), .B(_1070__bF_buf2), .C(regs_29__17_), .Y(_1088_) );
OAI21X1 OAI21X1_2213 ( .gnd(gnd), .vdd(vdd), .A(_1035__bF_buf2), .B(_1069__bF_buf2), .C(_1088_), .Y(_680_) );
OAI21X1 OAI21X1_2214 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf5), .B(_1070__bF_buf1), .C(regs_29__18_), .Y(_1089_) );
OAI21X1 OAI21X1_2215 ( .gnd(gnd), .vdd(vdd), .A(_1037__bF_buf2), .B(_1069__bF_buf1), .C(_1089_), .Y(_681_) );
OAI21X1 OAI21X1_2216 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_1070__bF_buf0), .C(regs_29__19_), .Y(_1090_) );
OAI21X1 OAI21X1_2217 ( .gnd(gnd), .vdd(vdd), .A(_1039__bF_buf2), .B(_1069__bF_buf0), .C(_1090_), .Y(_682_) );
OAI21X1 OAI21X1_2218 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf3), .B(_1070__bF_buf10), .C(regs_29__20_), .Y(_1091_) );
OAI21X1 OAI21X1_2219 ( .gnd(gnd), .vdd(vdd), .A(_1041__bF_buf2), .B(_1069__bF_buf4), .C(_1091_), .Y(_684_) );
OAI21X1 OAI21X1_2220 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf2), .B(_1070__bF_buf9), .C(regs_29__21_), .Y(_1092_) );
OAI21X1 OAI21X1_2221 ( .gnd(gnd), .vdd(vdd), .A(_1043__bF_buf2), .B(_1069__bF_buf3), .C(_1092_), .Y(_685_) );
OAI21X1 OAI21X1_2222 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1070__bF_buf8), .C(regs_29__22_), .Y(_1093_) );
OAI21X1 OAI21X1_2223 ( .gnd(gnd), .vdd(vdd), .A(_1045__bF_buf2), .B(_1069__bF_buf2), .C(_1093_), .Y(_686_) );
OAI21X1 OAI21X1_2224 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf0), .B(_1070__bF_buf7), .C(regs_29__23_), .Y(_1094_) );
OAI21X1 OAI21X1_2225 ( .gnd(gnd), .vdd(vdd), .A(_1047__bF_buf2), .B(_1069__bF_buf1), .C(_1094_), .Y(_687_) );
OAI21X1 OAI21X1_2226 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf7), .B(_1070__bF_buf6), .C(regs_29__24_), .Y(_1095_) );
OAI21X1 OAI21X1_2227 ( .gnd(gnd), .vdd(vdd), .A(_1049__bF_buf2), .B(_1069__bF_buf0), .C(_1095_), .Y(_688_) );
OAI21X1 OAI21X1_2228 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf6), .B(_1070__bF_buf5), .C(regs_29__25_), .Y(_1096_) );
OAI21X1 OAI21X1_2229 ( .gnd(gnd), .vdd(vdd), .A(_1051__bF_buf2), .B(_1069__bF_buf4), .C(_1096_), .Y(_689_) );
OAI21X1 OAI21X1_2230 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf5), .B(_1070__bF_buf4), .C(regs_29__26_), .Y(_1097_) );
OAI21X1 OAI21X1_2231 ( .gnd(gnd), .vdd(vdd), .A(_1053__bF_buf2), .B(_1069__bF_buf3), .C(_1097_), .Y(_690_) );
OAI21X1 OAI21X1_2232 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf4), .B(_1070__bF_buf3), .C(regs_29__27_), .Y(_1098_) );
OAI21X1 OAI21X1_2233 ( .gnd(gnd), .vdd(vdd), .A(_1055__bF_buf2), .B(_1069__bF_buf2), .C(_1098_), .Y(_691_) );
OAI21X1 OAI21X1_2234 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf3), .B(_1070__bF_buf2), .C(regs_29__28_), .Y(_1099_) );
OAI21X1 OAI21X1_2235 ( .gnd(gnd), .vdd(vdd), .A(_1057__bF_buf2), .B(_1069__bF_buf1), .C(_1099_), .Y(_692_) );
OAI21X1 OAI21X1_2236 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf2), .B(_1070__bF_buf1), .C(regs_29__29_), .Y(_1100_) );
OAI21X1 OAI21X1_2237 ( .gnd(gnd), .vdd(vdd), .A(_1059__bF_buf2), .B(_1069__bF_buf0), .C(_1100_), .Y(_693_) );
OAI21X1 OAI21X1_2238 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf1), .B(_1070__bF_buf0), .C(regs_29__30_), .Y(_1101_) );
OAI21X1 OAI21X1_2239 ( .gnd(gnd), .vdd(vdd), .A(_1061__bF_buf2), .B(_1069__bF_buf4), .C(_1101_), .Y(_695_) );
OAI21X1 OAI21X1_2240 ( .gnd(gnd), .vdd(vdd), .A(_1000__bF_buf0), .B(_1070__bF_buf10), .C(regs_29__31_), .Y(_1102_) );
OAI21X1 OAI21X1_2241 ( .gnd(gnd), .vdd(vdd), .A(_1063__bF_buf2), .B(_1069__bF_buf3), .C(_1102_), .Y(_696_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(waddr[1]), .Y(_1103_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_997_), .B(_1103_), .Y(_1104_) );
NOR2X1 NOR2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf0), .B(_1000__bF_buf7), .Y(_1105_) );
NOR2X1 NOR2X1_251 ( .gnd(gnd), .vdd(vdd), .A(regs_28__0_), .B(_1105__bF_buf7), .Y(_1106_) );
AOI21X1 AOI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_992__bF_buf2), .B(_1105__bF_buf6), .C(_1106_), .Y(_640_) );
NOR2X1 NOR2X1_252 ( .gnd(gnd), .vdd(vdd), .A(regs_28__1_), .B(_1105__bF_buf5), .Y(_1107_) );
AOI21X1 AOI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_1003__bF_buf2), .B(_1105__bF_buf4), .C(_1107_), .Y(_651_) );
NOR2X1 NOR2X1_253 ( .gnd(gnd), .vdd(vdd), .A(regs_28__2_), .B(_1105__bF_buf3), .Y(_1108_) );
AOI21X1 AOI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf2), .B(_1105__bF_buf2), .C(_1108_), .Y(_662_) );
NOR2X1 NOR2X1_254 ( .gnd(gnd), .vdd(vdd), .A(regs_28__3_), .B(_1105__bF_buf1), .Y(_1109_) );
AOI21X1 AOI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_1007__bF_buf2), .B(_1105__bF_buf0), .C(_1109_), .Y(_665_) );
NOR2X1 NOR2X1_255 ( .gnd(gnd), .vdd(vdd), .A(regs_28__4_), .B(_1105__bF_buf7), .Y(_1110_) );
AOI21X1 AOI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_1009__bF_buf1), .B(_1105__bF_buf6), .C(_1110_), .Y(_666_) );
NOR2X1 NOR2X1_256 ( .gnd(gnd), .vdd(vdd), .A(regs_28__5_), .B(_1105__bF_buf5), .Y(_1111_) );
AOI21X1 AOI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_1011__bF_buf1), .B(_1105__bF_buf4), .C(_1111_), .Y(_667_) );
NOR2X1 NOR2X1_257 ( .gnd(gnd), .vdd(vdd), .A(regs_28__6_), .B(_1105__bF_buf3), .Y(_1112_) );
AOI21X1 AOI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_1013__bF_buf1), .B(_1105__bF_buf2), .C(_1112_), .Y(_668_) );
NOR2X1 NOR2X1_258 ( .gnd(gnd), .vdd(vdd), .A(regs_28__7_), .B(_1105__bF_buf1), .Y(_1113_) );
AOI21X1 AOI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_1015__bF_buf1), .B(_1105__bF_buf0), .C(_1113_), .Y(_669_) );
NOR2X1 NOR2X1_259 ( .gnd(gnd), .vdd(vdd), .A(regs_28__8_), .B(_1105__bF_buf7), .Y(_1114_) );
AOI21X1 AOI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf1), .B(_1105__bF_buf6), .C(_1114_), .Y(_670_) );
NOR2X1 NOR2X1_260 ( .gnd(gnd), .vdd(vdd), .A(regs_28__9_), .B(_1105__bF_buf5), .Y(_1115_) );
AOI21X1 AOI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_1019__bF_buf1), .B(_1105__bF_buf4), .C(_1115_), .Y(_671_) );
NOR2X1 NOR2X1_261 ( .gnd(gnd), .vdd(vdd), .A(regs_28__10_), .B(_1105__bF_buf3), .Y(_1116_) );
AOI21X1 AOI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_1021__bF_buf1), .B(_1105__bF_buf2), .C(_1116_), .Y(_641_) );
NOR2X1 NOR2X1_262 ( .gnd(gnd), .vdd(vdd), .A(regs_28__11_), .B(_1105__bF_buf1), .Y(_1117_) );
AOI21X1 AOI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_1023__bF_buf1), .B(_1105__bF_buf0), .C(_1117_), .Y(_642_) );
NOR2X1 NOR2X1_263 ( .gnd(gnd), .vdd(vdd), .A(regs_28__12_), .B(_1105__bF_buf7), .Y(_1118_) );
AOI21X1 AOI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_1025__bF_buf1), .B(_1105__bF_buf6), .C(_1118_), .Y(_643_) );
NOR2X1 NOR2X1_264 ( .gnd(gnd), .vdd(vdd), .A(regs_28__13_), .B(_1105__bF_buf5), .Y(_1119_) );
AOI21X1 AOI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_1027__bF_buf1), .B(_1105__bF_buf4), .C(_1119_), .Y(_644_) );
NOR2X1 NOR2X1_265 ( .gnd(gnd), .vdd(vdd), .A(regs_28__14_), .B(_1105__bF_buf3), .Y(_1120_) );
AOI21X1 AOI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_1029__bF_buf1), .B(_1105__bF_buf2), .C(_1120_), .Y(_645_) );
NOR2X1 NOR2X1_266 ( .gnd(gnd), .vdd(vdd), .A(regs_28__15_), .B(_1105__bF_buf1), .Y(_1121_) );
AOI21X1 AOI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf1), .B(_1105__bF_buf0), .C(_1121_), .Y(_646_) );
NOR2X1 NOR2X1_267 ( .gnd(gnd), .vdd(vdd), .A(regs_28__16_), .B(_1105__bF_buf7), .Y(_1122_) );
AOI21X1 AOI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_1033__bF_buf1), .B(_1105__bF_buf6), .C(_1122_), .Y(_647_) );
NOR2X1 NOR2X1_268 ( .gnd(gnd), .vdd(vdd), .A(regs_28__17_), .B(_1105__bF_buf5), .Y(_1123_) );
AOI21X1 AOI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_1035__bF_buf1), .B(_1105__bF_buf4), .C(_1123_), .Y(_648_) );
NOR2X1 NOR2X1_269 ( .gnd(gnd), .vdd(vdd), .A(regs_28__18_), .B(_1105__bF_buf3), .Y(_1124_) );
AOI21X1 AOI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_1037__bF_buf1), .B(_1105__bF_buf2), .C(_1124_), .Y(_649_) );
NOR2X1 NOR2X1_270 ( .gnd(gnd), .vdd(vdd), .A(regs_28__19_), .B(_1105__bF_buf1), .Y(_1125_) );
AOI21X1 AOI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_1039__bF_buf1), .B(_1105__bF_buf0), .C(_1125_), .Y(_650_) );
NOR2X1 NOR2X1_271 ( .gnd(gnd), .vdd(vdd), .A(regs_28__20_), .B(_1105__bF_buf7), .Y(_1126_) );
AOI21X1 AOI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_1041__bF_buf1), .B(_1105__bF_buf6), .C(_1126_), .Y(_652_) );
NOR2X1 NOR2X1_272 ( .gnd(gnd), .vdd(vdd), .A(regs_28__21_), .B(_1105__bF_buf5), .Y(_1127_) );
AOI21X1 AOI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_1043__bF_buf1), .B(_1105__bF_buf4), .C(_1127_), .Y(_653_) );
NOR2X1 NOR2X1_273 ( .gnd(gnd), .vdd(vdd), .A(regs_28__22_), .B(_1105__bF_buf3), .Y(_1128_) );
AOI21X1 AOI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_1045__bF_buf1), .B(_1105__bF_buf2), .C(_1128_), .Y(_654_) );
NOR2X1 NOR2X1_274 ( .gnd(gnd), .vdd(vdd), .A(regs_28__23_), .B(_1105__bF_buf1), .Y(_1129_) );
AOI21X1 AOI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_1047__bF_buf1), .B(_1105__bF_buf0), .C(_1129_), .Y(_655_) );
NOR2X1 NOR2X1_275 ( .gnd(gnd), .vdd(vdd), .A(regs_28__24_), .B(_1105__bF_buf7), .Y(_1130_) );
AOI21X1 AOI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_1049__bF_buf1), .B(_1105__bF_buf6), .C(_1130_), .Y(_656_) );
NOR2X1 NOR2X1_276 ( .gnd(gnd), .vdd(vdd), .A(regs_28__25_), .B(_1105__bF_buf5), .Y(_1131_) );
AOI21X1 AOI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_1051__bF_buf1), .B(_1105__bF_buf4), .C(_1131_), .Y(_657_) );
NOR2X1 NOR2X1_277 ( .gnd(gnd), .vdd(vdd), .A(regs_28__26_), .B(_1105__bF_buf3), .Y(_1132_) );
AOI21X1 AOI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_1053__bF_buf1), .B(_1105__bF_buf2), .C(_1132_), .Y(_658_) );
NOR2X1 NOR2X1_278 ( .gnd(gnd), .vdd(vdd), .A(regs_28__27_), .B(_1105__bF_buf1), .Y(_1133_) );
AOI21X1 AOI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_1055__bF_buf1), .B(_1105__bF_buf0), .C(_1133_), .Y(_659_) );
NOR2X1 NOR2X1_279 ( .gnd(gnd), .vdd(vdd), .A(regs_28__28_), .B(_1105__bF_buf7), .Y(_1134_) );
AOI21X1 AOI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_1057__bF_buf1), .B(_1105__bF_buf6), .C(_1134_), .Y(_660_) );
NOR2X1 NOR2X1_280 ( .gnd(gnd), .vdd(vdd), .A(regs_28__29_), .B(_1105__bF_buf5), .Y(_1135_) );
AOI21X1 AOI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_1059__bF_buf1), .B(_1105__bF_buf4), .C(_1135_), .Y(_661_) );
NOR2X1 NOR2X1_281 ( .gnd(gnd), .vdd(vdd), .A(regs_28__30_), .B(_1105__bF_buf3), .Y(_1136_) );
AOI21X1 AOI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_1061__bF_buf1), .B(_1105__bF_buf2), .C(_1136_), .Y(_663_) );
NOR2X1 NOR2X1_282 ( .gnd(gnd), .vdd(vdd), .A(regs_28__31_), .B(_1105__bF_buf1), .Y(_1137_) );
AOI21X1 AOI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_1063__bF_buf1), .B(_1105__bF_buf0), .C(_1137_), .Y(_664_) );
INVX2 INVX2_289 ( .gnd(gnd), .vdd(vdd), .A(regs_27__0_), .Y(_1138_) );
INVX2 INVX2_290 ( .gnd(gnd), .vdd(vdd), .A(waddr[2]), .Y(_1139_) );
NOR2X1 NOR2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_1139_), .B(_995_), .Y(_1140_) );
INVX8 INVX8_43 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .Y(_1141_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(wen), .B(_1103_), .C(_1066_), .Y(_1142_) );
NOR2X1 NOR2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_1142__bF_buf3), .B(_1141__bF_buf3), .Y(_1143_) );
NAND2X1 NAND2X1_1105 ( .gnd(gnd), .vdd(vdd), .A(wdata[0]), .B(_1143__bF_buf7), .Y(_1144_) );
OAI21X1 OAI21X1_2242 ( .gnd(gnd), .vdd(vdd), .A(_1138_), .B(_1143__bF_buf6), .C(_1144_), .Y(_608_) );
INVX2 INVX2_291 ( .gnd(gnd), .vdd(vdd), .A(regs_27__1_), .Y(_1145_) );
NAND2X1 NAND2X1_1106 ( .gnd(gnd), .vdd(vdd), .A(wdata[1]), .B(_1143__bF_buf5), .Y(_1146_) );
OAI21X1 OAI21X1_2243 ( .gnd(gnd), .vdd(vdd), .A(_1145_), .B(_1143__bF_buf4), .C(_1146_), .Y(_619_) );
INVX2 INVX2_292 ( .gnd(gnd), .vdd(vdd), .A(regs_27__2_), .Y(_1147_) );
NAND2X1 NAND2X1_1107 ( .gnd(gnd), .vdd(vdd), .A(wdata[2]), .B(_1143__bF_buf3), .Y(_1148_) );
OAI21X1 OAI21X1_2244 ( .gnd(gnd), .vdd(vdd), .A(_1147_), .B(_1143__bF_buf2), .C(_1148_), .Y(_630_) );
INVX2 INVX2_293 ( .gnd(gnd), .vdd(vdd), .A(regs_27__3_), .Y(_1149_) );
NAND2X1 NAND2X1_1108 ( .gnd(gnd), .vdd(vdd), .A(wdata[3]), .B(_1143__bF_buf1), .Y(_1150_) );
OAI21X1 OAI21X1_2245 ( .gnd(gnd), .vdd(vdd), .A(_1149_), .B(_1143__bF_buf0), .C(_1150_), .Y(_633_) );
INVX2 INVX2_294 ( .gnd(gnd), .vdd(vdd), .A(regs_27__4_), .Y(_1151_) );
NAND2X1 NAND2X1_1109 ( .gnd(gnd), .vdd(vdd), .A(wdata[4]), .B(_1143__bF_buf7), .Y(_1152_) );
OAI21X1 OAI21X1_2246 ( .gnd(gnd), .vdd(vdd), .A(_1151_), .B(_1143__bF_buf6), .C(_1152_), .Y(_634_) );
INVX2 INVX2_295 ( .gnd(gnd), .vdd(vdd), .A(regs_27__5_), .Y(_1153_) );
NAND2X1 NAND2X1_1110 ( .gnd(gnd), .vdd(vdd), .A(wdata[5]), .B(_1143__bF_buf5), .Y(_1154_) );
OAI21X1 OAI21X1_2247 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(_1143__bF_buf4), .C(_1154_), .Y(_635_) );
INVX2 INVX2_296 ( .gnd(gnd), .vdd(vdd), .A(regs_27__6_), .Y(_1155_) );
NAND2X1 NAND2X1_1111 ( .gnd(gnd), .vdd(vdd), .A(wdata[6]), .B(_1143__bF_buf3), .Y(_1156_) );
OAI21X1 OAI21X1_2248 ( .gnd(gnd), .vdd(vdd), .A(_1155_), .B(_1143__bF_buf2), .C(_1156_), .Y(_636_) );
INVX2 INVX2_297 ( .gnd(gnd), .vdd(vdd), .A(regs_27__7_), .Y(_1157_) );
NAND2X1 NAND2X1_1112 ( .gnd(gnd), .vdd(vdd), .A(wdata[7]), .B(_1143__bF_buf1), .Y(_1158_) );
OAI21X1 OAI21X1_2249 ( .gnd(gnd), .vdd(vdd), .A(_1157_), .B(_1143__bF_buf0), .C(_1158_), .Y(_637_) );
INVX2 INVX2_298 ( .gnd(gnd), .vdd(vdd), .A(regs_27__8_), .Y(_1159_) );
NAND2X1 NAND2X1_1113 ( .gnd(gnd), .vdd(vdd), .A(wdata[8]), .B(_1143__bF_buf7), .Y(_1160_) );
OAI21X1 OAI21X1_2250 ( .gnd(gnd), .vdd(vdd), .A(_1159_), .B(_1143__bF_buf6), .C(_1160_), .Y(_638_) );
INVX2 INVX2_299 ( .gnd(gnd), .vdd(vdd), .A(regs_27__9_), .Y(_1161_) );
NAND2X1 NAND2X1_1114 ( .gnd(gnd), .vdd(vdd), .A(wdata[9]), .B(_1143__bF_buf5), .Y(_1162_) );
OAI21X1 OAI21X1_2251 ( .gnd(gnd), .vdd(vdd), .A(_1161_), .B(_1143__bF_buf4), .C(_1162_), .Y(_639_) );
INVX2 INVX2_300 ( .gnd(gnd), .vdd(vdd), .A(regs_27__10_), .Y(_1163_) );
NAND2X1 NAND2X1_1115 ( .gnd(gnd), .vdd(vdd), .A(wdata[10]), .B(_1143__bF_buf3), .Y(_1164_) );
OAI21X1 OAI21X1_2252 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(_1143__bF_buf2), .C(_1164_), .Y(_609_) );
INVX2 INVX2_301 ( .gnd(gnd), .vdd(vdd), .A(regs_27__11_), .Y(_1165_) );
NAND2X1 NAND2X1_1116 ( .gnd(gnd), .vdd(vdd), .A(wdata[11]), .B(_1143__bF_buf1), .Y(_1166_) );
OAI21X1 OAI21X1_2253 ( .gnd(gnd), .vdd(vdd), .A(_1165_), .B(_1143__bF_buf0), .C(_1166_), .Y(_610_) );
INVX2 INVX2_302 ( .gnd(gnd), .vdd(vdd), .A(regs_27__12_), .Y(_1167_) );
NAND2X1 NAND2X1_1117 ( .gnd(gnd), .vdd(vdd), .A(wdata[12]), .B(_1143__bF_buf7), .Y(_1168_) );
OAI21X1 OAI21X1_2254 ( .gnd(gnd), .vdd(vdd), .A(_1167_), .B(_1143__bF_buf6), .C(_1168_), .Y(_611_) );
INVX2 INVX2_303 ( .gnd(gnd), .vdd(vdd), .A(regs_27__13_), .Y(_1169_) );
NAND2X1 NAND2X1_1118 ( .gnd(gnd), .vdd(vdd), .A(wdata[13]), .B(_1143__bF_buf5), .Y(_1170_) );
OAI21X1 OAI21X1_2255 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_1143__bF_buf4), .C(_1170_), .Y(_612_) );
INVX2 INVX2_304 ( .gnd(gnd), .vdd(vdd), .A(regs_27__14_), .Y(_1171_) );
NAND2X1 NAND2X1_1119 ( .gnd(gnd), .vdd(vdd), .A(wdata[14]), .B(_1143__bF_buf3), .Y(_1172_) );
OAI21X1 OAI21X1_2256 ( .gnd(gnd), .vdd(vdd), .A(_1171_), .B(_1143__bF_buf2), .C(_1172_), .Y(_613_) );
INVX2 INVX2_305 ( .gnd(gnd), .vdd(vdd), .A(regs_27__15_), .Y(_1173_) );
NAND2X1 NAND2X1_1120 ( .gnd(gnd), .vdd(vdd), .A(wdata[15]), .B(_1143__bF_buf1), .Y(_1174_) );
OAI21X1 OAI21X1_2257 ( .gnd(gnd), .vdd(vdd), .A(_1173_), .B(_1143__bF_buf0), .C(_1174_), .Y(_614_) );
INVX2 INVX2_306 ( .gnd(gnd), .vdd(vdd), .A(regs_27__16_), .Y(_1175_) );
NAND2X1 NAND2X1_1121 ( .gnd(gnd), .vdd(vdd), .A(wdata[16]), .B(_1143__bF_buf7), .Y(_1176_) );
OAI21X1 OAI21X1_2258 ( .gnd(gnd), .vdd(vdd), .A(_1175_), .B(_1143__bF_buf6), .C(_1176_), .Y(_615_) );
INVX2 INVX2_307 ( .gnd(gnd), .vdd(vdd), .A(regs_27__17_), .Y(_1177_) );
NAND2X1 NAND2X1_1122 ( .gnd(gnd), .vdd(vdd), .A(wdata[17]), .B(_1143__bF_buf5), .Y(_1178_) );
OAI21X1 OAI21X1_2259 ( .gnd(gnd), .vdd(vdd), .A(_1177_), .B(_1143__bF_buf4), .C(_1178_), .Y(_616_) );
INVX2 INVX2_308 ( .gnd(gnd), .vdd(vdd), .A(regs_27__18_), .Y(_1179_) );
NAND2X1 NAND2X1_1123 ( .gnd(gnd), .vdd(vdd), .A(wdata[18]), .B(_1143__bF_buf3), .Y(_1180_) );
OAI21X1 OAI21X1_2260 ( .gnd(gnd), .vdd(vdd), .A(_1179_), .B(_1143__bF_buf2), .C(_1180_), .Y(_617_) );
INVX2 INVX2_309 ( .gnd(gnd), .vdd(vdd), .A(regs_27__19_), .Y(_1181_) );
NAND2X1 NAND2X1_1124 ( .gnd(gnd), .vdd(vdd), .A(wdata[19]), .B(_1143__bF_buf1), .Y(_1182_) );
OAI21X1 OAI21X1_2261 ( .gnd(gnd), .vdd(vdd), .A(_1181_), .B(_1143__bF_buf0), .C(_1182_), .Y(_618_) );
INVX2 INVX2_310 ( .gnd(gnd), .vdd(vdd), .A(regs_27__20_), .Y(_1183_) );
NAND2X1 NAND2X1_1125 ( .gnd(gnd), .vdd(vdd), .A(wdata[20]), .B(_1143__bF_buf7), .Y(_1184_) );
OAI21X1 OAI21X1_2262 ( .gnd(gnd), .vdd(vdd), .A(_1183_), .B(_1143__bF_buf6), .C(_1184_), .Y(_620_) );
INVX2 INVX2_311 ( .gnd(gnd), .vdd(vdd), .A(regs_27__21_), .Y(_1185_) );
NAND2X1 NAND2X1_1126 ( .gnd(gnd), .vdd(vdd), .A(wdata[21]), .B(_1143__bF_buf5), .Y(_1186_) );
OAI21X1 OAI21X1_2263 ( .gnd(gnd), .vdd(vdd), .A(_1185_), .B(_1143__bF_buf4), .C(_1186_), .Y(_621_) );
INVX2 INVX2_312 ( .gnd(gnd), .vdd(vdd), .A(regs_27__22_), .Y(_1187_) );
NAND2X1 NAND2X1_1127 ( .gnd(gnd), .vdd(vdd), .A(wdata[22]), .B(_1143__bF_buf3), .Y(_1188_) );
OAI21X1 OAI21X1_2264 ( .gnd(gnd), .vdd(vdd), .A(_1187_), .B(_1143__bF_buf2), .C(_1188_), .Y(_622_) );
INVX2 INVX2_313 ( .gnd(gnd), .vdd(vdd), .A(regs_27__23_), .Y(_1189_) );
NAND2X1 NAND2X1_1128 ( .gnd(gnd), .vdd(vdd), .A(wdata[23]), .B(_1143__bF_buf1), .Y(_1190_) );
OAI21X1 OAI21X1_2265 ( .gnd(gnd), .vdd(vdd), .A(_1189_), .B(_1143__bF_buf0), .C(_1190_), .Y(_623_) );
INVX2 INVX2_314 ( .gnd(gnd), .vdd(vdd), .A(regs_27__24_), .Y(_1191_) );
NAND2X1 NAND2X1_1129 ( .gnd(gnd), .vdd(vdd), .A(wdata[24]), .B(_1143__bF_buf7), .Y(_1192_) );
OAI21X1 OAI21X1_2266 ( .gnd(gnd), .vdd(vdd), .A(_1191_), .B(_1143__bF_buf6), .C(_1192_), .Y(_624_) );
INVX2 INVX2_315 ( .gnd(gnd), .vdd(vdd), .A(regs_27__25_), .Y(_1193_) );
NAND2X1 NAND2X1_1130 ( .gnd(gnd), .vdd(vdd), .A(wdata[25]), .B(_1143__bF_buf5), .Y(_1194_) );
OAI21X1 OAI21X1_2267 ( .gnd(gnd), .vdd(vdd), .A(_1193_), .B(_1143__bF_buf4), .C(_1194_), .Y(_625_) );
INVX2 INVX2_316 ( .gnd(gnd), .vdd(vdd), .A(regs_27__26_), .Y(_1195_) );
NAND2X1 NAND2X1_1131 ( .gnd(gnd), .vdd(vdd), .A(wdata[26]), .B(_1143__bF_buf3), .Y(_1196_) );
OAI21X1 OAI21X1_2268 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(_1143__bF_buf2), .C(_1196_), .Y(_626_) );
INVX2 INVX2_317 ( .gnd(gnd), .vdd(vdd), .A(regs_27__27_), .Y(_1197_) );
NAND2X1 NAND2X1_1132 ( .gnd(gnd), .vdd(vdd), .A(wdata[27]), .B(_1143__bF_buf1), .Y(_1198_) );
OAI21X1 OAI21X1_2269 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(_1143__bF_buf0), .C(_1198_), .Y(_627_) );
INVX2 INVX2_318 ( .gnd(gnd), .vdd(vdd), .A(regs_27__28_), .Y(_1199_) );
NAND2X1 NAND2X1_1133 ( .gnd(gnd), .vdd(vdd), .A(wdata[28]), .B(_1143__bF_buf7), .Y(_1200_) );
OAI21X1 OAI21X1_2270 ( .gnd(gnd), .vdd(vdd), .A(_1199_), .B(_1143__bF_buf6), .C(_1200_), .Y(_628_) );
INVX2 INVX2_319 ( .gnd(gnd), .vdd(vdd), .A(regs_27__29_), .Y(_1201_) );
NAND2X1 NAND2X1_1134 ( .gnd(gnd), .vdd(vdd), .A(wdata[29]), .B(_1143__bF_buf5), .Y(_1202_) );
OAI21X1 OAI21X1_2271 ( .gnd(gnd), .vdd(vdd), .A(_1201_), .B(_1143__bF_buf4), .C(_1202_), .Y(_629_) );
INVX2 INVX2_320 ( .gnd(gnd), .vdd(vdd), .A(regs_27__30_), .Y(_1203_) );
NAND2X1 NAND2X1_1135 ( .gnd(gnd), .vdd(vdd), .A(wdata[30]), .B(_1143__bF_buf3), .Y(_1204_) );
OAI21X1 OAI21X1_2272 ( .gnd(gnd), .vdd(vdd), .A(_1203_), .B(_1143__bF_buf2), .C(_1204_), .Y(_631_) );
INVX2 INVX2_321 ( .gnd(gnd), .vdd(vdd), .A(regs_27__31_), .Y(_1205_) );
NAND2X1 NAND2X1_1136 ( .gnd(gnd), .vdd(vdd), .A(wdata[31]), .B(_1143__bF_buf1), .Y(_1206_) );
OAI21X1 OAI21X1_2273 ( .gnd(gnd), .vdd(vdd), .A(_1205_), .B(_1143__bF_buf0), .C(_1206_), .Y(_632_) );
NOR2X1 NOR2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_1001__bF_buf9), .B(_1141__bF_buf2), .Y(_1207_) );
NOR2X1 NOR2X1_286 ( .gnd(gnd), .vdd(vdd), .A(regs_26__0_), .B(_1207__bF_buf7), .Y(_1208_) );
AOI21X1 AOI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_992__bF_buf1), .B(_1207__bF_buf6), .C(_1208_), .Y(_576_) );
NOR2X1 NOR2X1_287 ( .gnd(gnd), .vdd(vdd), .A(regs_26__1_), .B(_1207__bF_buf5), .Y(_1209_) );
AOI21X1 AOI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_1003__bF_buf1), .B(_1207__bF_buf4), .C(_1209_), .Y(_587_) );
NOR2X1 NOR2X1_288 ( .gnd(gnd), .vdd(vdd), .A(regs_26__2_), .B(_1207__bF_buf3), .Y(_1210_) );
AOI21X1 AOI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf1), .B(_1207__bF_buf2), .C(_1210_), .Y(_598_) );
NOR2X1 NOR2X1_289 ( .gnd(gnd), .vdd(vdd), .A(regs_26__3_), .B(_1207__bF_buf1), .Y(_1211_) );
AOI21X1 AOI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_1007__bF_buf1), .B(_1207__bF_buf0), .C(_1211_), .Y(_601_) );
NOR2X1 NOR2X1_290 ( .gnd(gnd), .vdd(vdd), .A(regs_26__4_), .B(_1207__bF_buf7), .Y(_1212_) );
AOI21X1 AOI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_1009__bF_buf0), .B(_1207__bF_buf6), .C(_1212_), .Y(_602_) );
NOR2X1 NOR2X1_291 ( .gnd(gnd), .vdd(vdd), .A(regs_26__5_), .B(_1207__bF_buf5), .Y(_1213_) );
AOI21X1 AOI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_1011__bF_buf0), .B(_1207__bF_buf4), .C(_1213_), .Y(_603_) );
NOR2X1 NOR2X1_292 ( .gnd(gnd), .vdd(vdd), .A(regs_26__6_), .B(_1207__bF_buf3), .Y(_1214_) );
AOI21X1 AOI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_1013__bF_buf0), .B(_1207__bF_buf2), .C(_1214_), .Y(_604_) );
NOR2X1 NOR2X1_293 ( .gnd(gnd), .vdd(vdd), .A(regs_26__7_), .B(_1207__bF_buf1), .Y(_1215_) );
AOI21X1 AOI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_1015__bF_buf0), .B(_1207__bF_buf0), .C(_1215_), .Y(_605_) );
NOR2X1 NOR2X1_294 ( .gnd(gnd), .vdd(vdd), .A(regs_26__8_), .B(_1207__bF_buf7), .Y(_1216_) );
AOI21X1 AOI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf0), .B(_1207__bF_buf6), .C(_1216_), .Y(_606_) );
NOR2X1 NOR2X1_295 ( .gnd(gnd), .vdd(vdd), .A(regs_26__9_), .B(_1207__bF_buf5), .Y(_1217_) );
AOI21X1 AOI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_1019__bF_buf0), .B(_1207__bF_buf4), .C(_1217_), .Y(_607_) );
NOR2X1 NOR2X1_296 ( .gnd(gnd), .vdd(vdd), .A(regs_26__10_), .B(_1207__bF_buf3), .Y(_1218_) );
AOI21X1 AOI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_1021__bF_buf0), .B(_1207__bF_buf2), .C(_1218_), .Y(_577_) );
NOR2X1 NOR2X1_297 ( .gnd(gnd), .vdd(vdd), .A(regs_26__11_), .B(_1207__bF_buf1), .Y(_1219_) );
AOI21X1 AOI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(_1023__bF_buf0), .B(_1207__bF_buf0), .C(_1219_), .Y(_578_) );
NOR2X1 NOR2X1_298 ( .gnd(gnd), .vdd(vdd), .A(regs_26__12_), .B(_1207__bF_buf7), .Y(_1220_) );
AOI21X1 AOI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_1025__bF_buf0), .B(_1207__bF_buf6), .C(_1220_), .Y(_579_) );
NOR2X1 NOR2X1_299 ( .gnd(gnd), .vdd(vdd), .A(regs_26__13_), .B(_1207__bF_buf5), .Y(_1221_) );
AOI21X1 AOI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_1027__bF_buf0), .B(_1207__bF_buf4), .C(_1221_), .Y(_580_) );
NOR2X1 NOR2X1_300 ( .gnd(gnd), .vdd(vdd), .A(regs_26__14_), .B(_1207__bF_buf3), .Y(_1222_) );
AOI21X1 AOI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(_1029__bF_buf0), .B(_1207__bF_buf2), .C(_1222_), .Y(_581_) );
NOR2X1 NOR2X1_301 ( .gnd(gnd), .vdd(vdd), .A(regs_26__15_), .B(_1207__bF_buf1), .Y(_1223_) );
AOI21X1 AOI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf0), .B(_1207__bF_buf0), .C(_1223_), .Y(_582_) );
NOR2X1 NOR2X1_302 ( .gnd(gnd), .vdd(vdd), .A(regs_26__16_), .B(_1207__bF_buf7), .Y(_1224_) );
AOI21X1 AOI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_1033__bF_buf0), .B(_1207__bF_buf6), .C(_1224_), .Y(_583_) );
NOR2X1 NOR2X1_303 ( .gnd(gnd), .vdd(vdd), .A(regs_26__17_), .B(_1207__bF_buf5), .Y(_1225_) );
AOI21X1 AOI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_1035__bF_buf0), .B(_1207__bF_buf4), .C(_1225_), .Y(_584_) );
NOR2X1 NOR2X1_304 ( .gnd(gnd), .vdd(vdd), .A(regs_26__18_), .B(_1207__bF_buf3), .Y(_1226_) );
AOI21X1 AOI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_1037__bF_buf0), .B(_1207__bF_buf2), .C(_1226_), .Y(_585_) );
NOR2X1 NOR2X1_305 ( .gnd(gnd), .vdd(vdd), .A(regs_26__19_), .B(_1207__bF_buf1), .Y(_1227_) );
AOI21X1 AOI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_1039__bF_buf0), .B(_1207__bF_buf0), .C(_1227_), .Y(_586_) );
NOR2X1 NOR2X1_306 ( .gnd(gnd), .vdd(vdd), .A(regs_26__20_), .B(_1207__bF_buf7), .Y(_1228_) );
AOI21X1 AOI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_1041__bF_buf0), .B(_1207__bF_buf6), .C(_1228_), .Y(_588_) );
NOR2X1 NOR2X1_307 ( .gnd(gnd), .vdd(vdd), .A(regs_26__21_), .B(_1207__bF_buf5), .Y(_1229_) );
AOI21X1 AOI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_1043__bF_buf0), .B(_1207__bF_buf4), .C(_1229_), .Y(_589_) );
NOR2X1 NOR2X1_308 ( .gnd(gnd), .vdd(vdd), .A(regs_26__22_), .B(_1207__bF_buf3), .Y(_1230_) );
AOI21X1 AOI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_1045__bF_buf0), .B(_1207__bF_buf2), .C(_1230_), .Y(_590_) );
NOR2X1 NOR2X1_309 ( .gnd(gnd), .vdd(vdd), .A(regs_26__23_), .B(_1207__bF_buf1), .Y(_1231_) );
AOI21X1 AOI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_1047__bF_buf0), .B(_1207__bF_buf0), .C(_1231_), .Y(_591_) );
NOR2X1 NOR2X1_310 ( .gnd(gnd), .vdd(vdd), .A(regs_26__24_), .B(_1207__bF_buf7), .Y(_1232_) );
AOI21X1 AOI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_1049__bF_buf0), .B(_1207__bF_buf6), .C(_1232_), .Y(_592_) );
NOR2X1 NOR2X1_311 ( .gnd(gnd), .vdd(vdd), .A(regs_26__25_), .B(_1207__bF_buf5), .Y(_1233_) );
AOI21X1 AOI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_1051__bF_buf0), .B(_1207__bF_buf4), .C(_1233_), .Y(_593_) );
NOR2X1 NOR2X1_312 ( .gnd(gnd), .vdd(vdd), .A(regs_26__26_), .B(_1207__bF_buf3), .Y(_1234_) );
AOI21X1 AOI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_1053__bF_buf0), .B(_1207__bF_buf2), .C(_1234_), .Y(_594_) );
NOR2X1 NOR2X1_313 ( .gnd(gnd), .vdd(vdd), .A(regs_26__27_), .B(_1207__bF_buf1), .Y(_1235_) );
AOI21X1 AOI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_1055__bF_buf0), .B(_1207__bF_buf0), .C(_1235_), .Y(_595_) );
NOR2X1 NOR2X1_314 ( .gnd(gnd), .vdd(vdd), .A(regs_26__28_), .B(_1207__bF_buf7), .Y(_1236_) );
AOI21X1 AOI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_1057__bF_buf0), .B(_1207__bF_buf6), .C(_1236_), .Y(_596_) );
NOR2X1 NOR2X1_315 ( .gnd(gnd), .vdd(vdd), .A(regs_26__29_), .B(_1207__bF_buf5), .Y(_1237_) );
AOI21X1 AOI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_1059__bF_buf0), .B(_1207__bF_buf4), .C(_1237_), .Y(_597_) );
NOR2X1 NOR2X1_316 ( .gnd(gnd), .vdd(vdd), .A(regs_26__30_), .B(_1207__bF_buf3), .Y(_1238_) );
AOI21X1 AOI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_1061__bF_buf0), .B(_1207__bF_buf2), .C(_1238_), .Y(_599_) );
NOR2X1 NOR2X1_317 ( .gnd(gnd), .vdd(vdd), .A(regs_26__31_), .B(_1207__bF_buf1), .Y(_1239_) );
AOI21X1 AOI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_1063__bF_buf0), .B(_1207__bF_buf0), .C(_1239_), .Y(_600_) );
NAND2X1 NAND2X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_1140_), .Y(_1240_) );
OAI21X1 OAI21X1_2274 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf1), .B(_1070__bF_buf9), .C(regs_25__0_), .Y(_1241_) );
OAI21X1 OAI21X1_2275 ( .gnd(gnd), .vdd(vdd), .A(_992__bF_buf0), .B(_1240__bF_buf4), .C(_1241_), .Y(_544_) );
OAI21X1 OAI21X1_2276 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf0), .B(_1070__bF_buf8), .C(regs_25__1_), .Y(_1242_) );
OAI21X1 OAI21X1_2277 ( .gnd(gnd), .vdd(vdd), .A(_1003__bF_buf0), .B(_1240__bF_buf3), .C(_1242_), .Y(_555_) );
OAI21X1 OAI21X1_2278 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf7), .B(_1070__bF_buf7), .C(regs_25__2_), .Y(_1243_) );
OAI21X1 OAI21X1_2279 ( .gnd(gnd), .vdd(vdd), .A(_1005__bF_buf0), .B(_1240__bF_buf2), .C(_1243_), .Y(_566_) );
OAI21X1 OAI21X1_2280 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf6), .B(_1070__bF_buf6), .C(regs_25__3_), .Y(_1244_) );
OAI21X1 OAI21X1_2281 ( .gnd(gnd), .vdd(vdd), .A(_1007__bF_buf0), .B(_1240__bF_buf1), .C(_1244_), .Y(_569_) );
OAI21X1 OAI21X1_2282 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf5), .B(_1070__bF_buf5), .C(regs_25__4_), .Y(_1245_) );
OAI21X1 OAI21X1_2283 ( .gnd(gnd), .vdd(vdd), .A(_1009__bF_buf3), .B(_1240__bF_buf0), .C(_1245_), .Y(_570_) );
OAI21X1 OAI21X1_2284 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf4), .B(_1070__bF_buf4), .C(regs_25__5_), .Y(_1246_) );
OAI21X1 OAI21X1_2285 ( .gnd(gnd), .vdd(vdd), .A(_1011__bF_buf3), .B(_1240__bF_buf4), .C(_1246_), .Y(_571_) );
OAI21X1 OAI21X1_2286 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf3), .B(_1070__bF_buf3), .C(regs_25__6_), .Y(_1247_) );
OAI21X1 OAI21X1_2287 ( .gnd(gnd), .vdd(vdd), .A(_1013__bF_buf3), .B(_1240__bF_buf3), .C(_1247_), .Y(_572_) );
OAI21X1 OAI21X1_2288 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf2), .B(_1070__bF_buf2), .C(regs_25__7_), .Y(_1248_) );
OAI21X1 OAI21X1_2289 ( .gnd(gnd), .vdd(vdd), .A(_1015__bF_buf3), .B(_1240__bF_buf2), .C(_1248_), .Y(_573_) );
OAI21X1 OAI21X1_2290 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf1), .B(_1070__bF_buf1), .C(regs_25__8_), .Y(_1249_) );
OAI21X1 OAI21X1_2291 ( .gnd(gnd), .vdd(vdd), .A(_1017__bF_buf3), .B(_1240__bF_buf1), .C(_1249_), .Y(_574_) );
OAI21X1 OAI21X1_2292 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf0), .B(_1070__bF_buf0), .C(regs_25__9_), .Y(_1250_) );
OAI21X1 OAI21X1_2293 ( .gnd(gnd), .vdd(vdd), .A(_1019__bF_buf3), .B(_1240__bF_buf0), .C(_1250_), .Y(_575_) );
OAI21X1 OAI21X1_2294 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf7), .B(_1070__bF_buf10), .C(regs_25__10_), .Y(_1251_) );
OAI21X1 OAI21X1_2295 ( .gnd(gnd), .vdd(vdd), .A(_1021__bF_buf3), .B(_1240__bF_buf4), .C(_1251_), .Y(_545_) );
OAI21X1 OAI21X1_2296 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf6), .B(_1070__bF_buf9), .C(regs_25__11_), .Y(_1252_) );
OAI21X1 OAI21X1_2297 ( .gnd(gnd), .vdd(vdd), .A(_1023__bF_buf3), .B(_1240__bF_buf3), .C(_1252_), .Y(_546_) );
OAI21X1 OAI21X1_2298 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf5), .B(_1070__bF_buf8), .C(regs_25__12_), .Y(_1253_) );
OAI21X1 OAI21X1_2299 ( .gnd(gnd), .vdd(vdd), .A(_1025__bF_buf3), .B(_1240__bF_buf2), .C(_1253_), .Y(_547_) );
OAI21X1 OAI21X1_2300 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf4), .B(_1070__bF_buf7), .C(regs_25__13_), .Y(_1254_) );
OAI21X1 OAI21X1_2301 ( .gnd(gnd), .vdd(vdd), .A(_1027__bF_buf3), .B(_1240__bF_buf1), .C(_1254_), .Y(_548_) );
OAI21X1 OAI21X1_2302 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf3), .B(_1070__bF_buf6), .C(regs_25__14_), .Y(_1255_) );
OAI21X1 OAI21X1_2303 ( .gnd(gnd), .vdd(vdd), .A(_1029__bF_buf3), .B(_1240__bF_buf0), .C(_1255_), .Y(_549_) );
OAI21X1 OAI21X1_2304 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf2), .B(_1070__bF_buf5), .C(regs_25__15_), .Y(_1256_) );
OAI21X1 OAI21X1_2305 ( .gnd(gnd), .vdd(vdd), .A(_1031__bF_buf3), .B(_1240__bF_buf4), .C(_1256_), .Y(_550_) );
OAI21X1 OAI21X1_2306 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf1), .B(_1070__bF_buf4), .C(regs_25__16_), .Y(_1257_) );
OAI21X1 OAI21X1_2307 ( .gnd(gnd), .vdd(vdd), .A(_1033__bF_buf3), .B(_1240__bF_buf3), .C(_1257_), .Y(_551_) );
OAI21X1 OAI21X1_2308 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf0), .B(_1070__bF_buf3), .C(regs_25__17_), .Y(_1258_) );
OAI21X1 OAI21X1_2309 ( .gnd(gnd), .vdd(vdd), .A(_1035__bF_buf3), .B(_1240__bF_buf2), .C(_1258_), .Y(_552_) );
OAI21X1 OAI21X1_2310 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf7), .B(_1070__bF_buf2), .C(regs_25__18_), .Y(_1259_) );
OAI21X1 OAI21X1_2311 ( .gnd(gnd), .vdd(vdd), .A(_1037__bF_buf3), .B(_1240__bF_buf1), .C(_1259_), .Y(_553_) );
OAI21X1 OAI21X1_2312 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf6), .B(_1070__bF_buf1), .C(regs_25__19_), .Y(_1260_) );
OAI21X1 OAI21X1_2313 ( .gnd(gnd), .vdd(vdd), .A(_1039__bF_buf3), .B(_1240__bF_buf0), .C(_1260_), .Y(_554_) );
OAI21X1 OAI21X1_2314 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf5), .B(_1070__bF_buf0), .C(regs_25__20_), .Y(_1261_) );
OAI21X1 OAI21X1_2315 ( .gnd(gnd), .vdd(vdd), .A(_1041__bF_buf3), .B(_1240__bF_buf4), .C(_1261_), .Y(_556_) );
OAI21X1 OAI21X1_2316 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf4), .B(_1070__bF_buf10), .C(regs_25__21_), .Y(_1262_) );
OAI21X1 OAI21X1_2317 ( .gnd(gnd), .vdd(vdd), .A(_1043__bF_buf3), .B(_1240__bF_buf3), .C(_1262_), .Y(_557_) );
OAI21X1 OAI21X1_2318 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf3), .B(_1070__bF_buf9), .C(regs_25__22_), .Y(_1263_) );
OAI21X1 OAI21X1_2319 ( .gnd(gnd), .vdd(vdd), .A(_1045__bF_buf3), .B(_1240__bF_buf2), .C(_1263_), .Y(_558_) );
OAI21X1 OAI21X1_2320 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf2), .B(_1070__bF_buf8), .C(regs_25__23_), .Y(_1264_) );
OAI21X1 OAI21X1_2321 ( .gnd(gnd), .vdd(vdd), .A(_1047__bF_buf3), .B(_1240__bF_buf1), .C(_1264_), .Y(_559_) );
OAI21X1 OAI21X1_2322 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf1), .B(_1070__bF_buf7), .C(regs_25__24_), .Y(_1265_) );
OAI21X1 OAI21X1_2323 ( .gnd(gnd), .vdd(vdd), .A(_1049__bF_buf3), .B(_1240__bF_buf0), .C(_1265_), .Y(_560_) );
OAI21X1 OAI21X1_2324 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf0), .B(_1070__bF_buf6), .C(regs_25__25_), .Y(_1266_) );
OAI21X1 OAI21X1_2325 ( .gnd(gnd), .vdd(vdd), .A(_1051__bF_buf3), .B(_1240__bF_buf4), .C(_1266_), .Y(_561_) );
OAI21X1 OAI21X1_2326 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf7), .B(_1070__bF_buf5), .C(regs_25__26_), .Y(_1267_) );
OAI21X1 OAI21X1_2327 ( .gnd(gnd), .vdd(vdd), .A(_1053__bF_buf3), .B(_1240__bF_buf3), .C(_1267_), .Y(_562_) );
OAI21X1 OAI21X1_2328 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf6), .B(_1070__bF_buf4), .C(regs_25__27_), .Y(_1268_) );
OAI21X1 OAI21X1_2329 ( .gnd(gnd), .vdd(vdd), .A(_1055__bF_buf3), .B(_1240__bF_buf2), .C(_1268_), .Y(_563_) );
OAI21X1 OAI21X1_2330 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf5), .B(_1070__bF_buf3), .C(regs_25__28_), .Y(_1269_) );
OAI21X1 OAI21X1_2331 ( .gnd(gnd), .vdd(vdd), .A(_1057__bF_buf3), .B(_1240__bF_buf1), .C(_1269_), .Y(_564_) );
OAI21X1 OAI21X1_2332 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf4), .B(_1070__bF_buf2), .C(regs_25__29_), .Y(_1270_) );
OAI21X1 OAI21X1_2333 ( .gnd(gnd), .vdd(vdd), .A(_1059__bF_buf3), .B(_1240__bF_buf0), .C(_1270_), .Y(_565_) );
OAI21X1 OAI21X1_2334 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf3), .B(_1070__bF_buf1), .C(regs_25__30_), .Y(_1271_) );
OAI21X1 OAI21X1_2335 ( .gnd(gnd), .vdd(vdd), .A(_1061__bF_buf3), .B(_1240__bF_buf4), .C(_1271_), .Y(_567_) );
OAI21X1 OAI21X1_2336 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf2), .B(_1070__bF_buf0), .C(regs_25__31_), .Y(_1272_) );
OAI21X1 OAI21X1_2337 ( .gnd(gnd), .vdd(vdd), .A(_1063__bF_buf3), .B(_1240__bF_buf3), .C(_1272_), .Y(_568_) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(_1104__bF_buf14), .Y(_1273_) );
NAND2X1 NAND2X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_1273_), .Y(_1274_) );
OAI21X1 OAI21X1_2338 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf1), .B(_1104__bF_buf13), .C(regs_24__0_), .Y(_1275_) );
OAI21X1 OAI21X1_2339 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf1), .B(_992__bF_buf3), .C(_1275_), .Y(_512_) );
OAI21X1 OAI21X1_2340 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf0), .B(_1104__bF_buf12), .C(regs_24__1_), .Y(_1276_) );
OAI21X1 OAI21X1_2341 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf0), .B(_1003__bF_buf3), .C(_1276_), .Y(_523_) );
OAI21X1 OAI21X1_2342 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf7), .B(_1104__bF_buf11), .C(regs_24__2_), .Y(_1277_) );
OAI21X1 OAI21X1_2343 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf4), .B(_1005__bF_buf3), .C(_1277_), .Y(_534_) );
OAI21X1 OAI21X1_2344 ( .gnd(gnd), .vdd(vdd), .A(_1141__bF_buf6), .B(_1104__bF_buf10), .C(regs_24__3_), .Y(_1278_) );
OAI21X1 OAI21X1_2345 ( .gnd(gnd), .vdd(vdd), .A(_1274__bF_buf3), .B(_1007__bF_buf3), .C(_1278_), .Y(_537_) );
endmodule
