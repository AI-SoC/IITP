module add ( gnd, vdd, a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, rst, on, clk, out);

input gnd, vdd;
input a;
input b;
input c;
input d;
input e;
input f;
input g;
input h;
input i;
input j;
input k;
input l;
input m;
input n;
input o;
input p;
input q;
input r;
input s;
input t;
input u;
input v;
input w;
input x;
input y;
input z;
input rst;
input on;
input clk;
output out;

CLKBUF1 CLKBUF1_1 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf3) );
CLKBUF1 CLKBUF1_2 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf2) );
CLKBUF1 CLKBUF1_3 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf1) );
CLKBUF1 CLKBUF1_4 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf0) );
BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(_49_), .Y(_49__bF_buf5) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(_49_), .Y(_49__bF_buf4) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(_49_), .Y(_49__bF_buf3) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(_49_), .Y(_49__bF_buf2) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(_49_), .Y(_49__bF_buf1) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(_49_), .Y(_49__bF_buf0) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_49__bF_buf5), .C(_23_), .Y(_15_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(b1), .B(q), .Y(_24_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(b2), .B(_49__bF_buf4), .Y(_25_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_49__bF_buf3), .C(_25_), .Y(_14_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(k), .B(a8), .Y(_26_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(a9), .B(_49__bF_buf2), .Y(_27_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_49__bF_buf1), .C(_27_), .Y(_10_) );
XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(m), .B(a10), .Y(_28_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(a11), .B(_49__bF_buf0), .Y(_29_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_49__bF_buf5), .C(_29_), .Y(_1_) );
XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(a9), .B(l), .Y(_30_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(a10), .B(_49__bF_buf4), .Y(_31_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_49__bF_buf3), .C(_31_), .Y(_0_) );
XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(g), .B(a5), .Y(_32_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(a6), .B(_49__bF_buf2), .Y(_33_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_49__bF_buf1), .C(_33_), .Y(_7_) );
XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(j), .B(a7), .Y(_34_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(a8), .B(_49__bF_buf0), .Y(_35_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_49__bF_buf5), .C(_35_), .Y(_9_) );
XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(a6), .B(h), .Y(_36_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(a7), .B(_49__bF_buf4), .Y(_37_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_49__bF_buf3), .C(_37_), .Y(_8_) );
XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(d), .B(a2), .Y(_38_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(a3), .B(_49__bF_buf2), .Y(_39_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_49__bF_buf1), .C(_39_), .Y(_4_) );
XNOR2X1 XNOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(f), .B(a4), .Y(_40_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(a5), .B(_49__bF_buf0), .Y(_41_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_49__bF_buf5), .C(_41_), .Y(_6_) );
XNOR2X1 XNOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(a3), .B(e), .Y(_42_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(a4), .B(_49__bF_buf4), .Y(_43_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_49__bF_buf3), .C(_43_), .Y(_5_) );
XNOR2X1 XNOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(c), .B(a1), .Y(_44_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(a2), .B(_49__bF_buf2), .Y(_45_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_49__bF_buf1), .C(_45_), .Y(_3_) );
XNOR2X1 XNOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(a), .B(b), .Y(_46_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(a1), .B(_49__bF_buf0), .Y(_47_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_49__bF_buf5), .C(_47_), .Y(_2_) );
XNOR2X1 XNOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(b11), .B(a11), .Y(_48_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_49__bF_buf4), .B(_48_), .Y(_22_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_69_), .Y(out) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_22_), .Q(_69_) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_2_), .Q(a1) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3_), .Q(a2) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_4_), .Q(a3) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_5_), .Q(a4) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_6_), .Q(a5) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_7_), .Q(a6) );
DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_8_), .Q(a7) );
DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_9_), .Q(a8) );
DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_10_), .Q(a9) );
DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0_), .Q(a10) );
DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_1_), .Q(a11) );
DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_13_), .Q(b1) );
DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_14_), .Q(b2) );
DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_15_), .Q(b3) );
DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_16_), .Q(b4) );
DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_17_), .Q(b5) );
DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_18_), .Q(b6) );
DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_19_), .Q(b7) );
DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_20_), .Q(b8) );
DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_21_), .Q(b9) );
DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_11_), .Q(b10) );
DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_12_), .Q(b11) );
INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(_49_) );
XNOR2X1 XNOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(z), .B(b10), .Y(_50_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(b11), .B(_49__bF_buf3), .Y(_51_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_49__bF_buf2), .C(_51_), .Y(_12_) );
XNOR2X1 XNOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(y), .B(b9), .Y(_52_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(b10), .B(_49__bF_buf1), .Y(_53_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_49__bF_buf0), .C(_53_), .Y(_11_) );
XNOR2X1 XNOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(v), .B(b6), .Y(_54_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(b7), .B(_49__bF_buf5), .Y(_55_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_49__bF_buf4), .C(_55_), .Y(_19_) );
XNOR2X1 XNOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(x), .B(b8), .Y(_56_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(b9), .B(_49__bF_buf3), .Y(_57_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_49__bF_buf2), .C(_57_), .Y(_21_) );
XNOR2X1 XNOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(b7), .B(w), .Y(_58_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(b8), .B(_49__bF_buf1), .Y(_59_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_49__bF_buf0), .C(_59_), .Y(_20_) );
XNOR2X1 XNOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(s), .B(b3), .Y(_60_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(b4), .B(_49__bF_buf5), .Y(_61_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_49__bF_buf4), .C(_61_), .Y(_16_) );
XNOR2X1 XNOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(u), .B(b5), .Y(_62_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(b6), .B(_49__bF_buf3), .Y(_63_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_49__bF_buf2), .C(_63_), .Y(_18_) );
XNOR2X1 XNOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(b4), .B(t), .Y(_64_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(b5), .B(_49__bF_buf1), .Y(_65_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_49__bF_buf0), .C(_65_), .Y(_17_) );
XNOR2X1 XNOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(n), .B(o), .Y(_66_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(b1), .B(_49__bF_buf5), .Y(_67_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_66_), .B(_49__bF_buf4), .C(_67_), .Y(_13_) );
XNOR2X1 XNOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(r), .B(b2), .Y(_68_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(b3), .B(_49__bF_buf3), .Y(_23_) );
endmodule
